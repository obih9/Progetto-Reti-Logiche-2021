
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

signal RAM: ram_type := (
			0 => std_logic_vector(to_unsigned( 128,8)),
			1 => std_logic_vector(to_unsigned( 128,8)),
			2 => std_logic_vector(to_unsigned( 18,8)),
			3 => std_logic_vector(to_unsigned( 61,8)),
			4 => std_logic_vector(to_unsigned( 91,8)),
			5 => std_logic_vector(to_unsigned( 219,8)),
			6 => std_logic_vector(to_unsigned( 130,8)),
			7 => std_logic_vector(to_unsigned( 91,8)),
			8 => std_logic_vector(to_unsigned( 50,8)),
			9 => std_logic_vector(to_unsigned( 128,8)),
			10 => std_logic_vector(to_unsigned( 189,8)),
			11 => std_logic_vector(to_unsigned( 200,8)),
			12 => std_logic_vector(to_unsigned( 184,8)),
			13 => std_logic_vector(to_unsigned( 39,8)),
			14 => std_logic_vector(to_unsigned( 56,8)),
			15 => std_logic_vector(to_unsigned( 16,8)),
			16 => std_logic_vector(to_unsigned( 174,8)),
			17 => std_logic_vector(to_unsigned( 144,8)),
			18 => std_logic_vector(to_unsigned( 1,8)),
			19 => std_logic_vector(to_unsigned( 29,8)),
			20 => std_logic_vector(to_unsigned( 207,8)),
			21 => std_logic_vector(to_unsigned( 51,8)),
			22 => std_logic_vector(to_unsigned( 212,8)),
			23 => std_logic_vector(to_unsigned( 126,8)),
			24 => std_logic_vector(to_unsigned( 201,8)),
			25 => std_logic_vector(to_unsigned( 183,8)),
			26 => std_logic_vector(to_unsigned( 232,8)),
			27 => std_logic_vector(to_unsigned( 223,8)),
			28 => std_logic_vector(to_unsigned( 205,8)),
			29 => std_logic_vector(to_unsigned( 39,8)),
			30 => std_logic_vector(to_unsigned( 198,8)),
			31 => std_logic_vector(to_unsigned( 167,8)),
			32 => std_logic_vector(to_unsigned( 19,8)),
			33 => std_logic_vector(to_unsigned( 200,8)),
			34 => std_logic_vector(to_unsigned( 64,8)),
			35 => std_logic_vector(to_unsigned( 30,8)),
			36 => std_logic_vector(to_unsigned( 93,8)),
			37 => std_logic_vector(to_unsigned( 90,8)),
			38 => std_logic_vector(to_unsigned( 168,8)),
			39 => std_logic_vector(to_unsigned( 144,8)),
			40 => std_logic_vector(to_unsigned( 110,8)),
			41 => std_logic_vector(to_unsigned( 152,8)),
			42 => std_logic_vector(to_unsigned( 221,8)),
			43 => std_logic_vector(to_unsigned( 78,8)),
			44 => std_logic_vector(to_unsigned( 103,8)),
			45 => std_logic_vector(to_unsigned( 190,8)),
			46 => std_logic_vector(to_unsigned( 76,8)),
			47 => std_logic_vector(to_unsigned( 203,8)),
			48 => std_logic_vector(to_unsigned( 209,8)),
			49 => std_logic_vector(to_unsigned( 9,8)),
			50 => std_logic_vector(to_unsigned( 7,8)),
			51 => std_logic_vector(to_unsigned( 1,8)),
			52 => std_logic_vector(to_unsigned( 146,8)),
			53 => std_logic_vector(to_unsigned( 255,8)),
			54 => std_logic_vector(to_unsigned( 145,8)),
			55 => std_logic_vector(to_unsigned( 51,8)),
			56 => std_logic_vector(to_unsigned( 35,8)),
			57 => std_logic_vector(to_unsigned( 97,8)),
			58 => std_logic_vector(to_unsigned( 120,8)),
			59 => std_logic_vector(to_unsigned( 88,8)),
			60 => std_logic_vector(to_unsigned( 48,8)),
			61 => std_logic_vector(to_unsigned( 91,8)),
			62 => std_logic_vector(to_unsigned( 207,8)),
			63 => std_logic_vector(to_unsigned( 200,8)),
			64 => std_logic_vector(to_unsigned( 195,8)),
			65 => std_logic_vector(to_unsigned( 69,8)),
			66 => std_logic_vector(to_unsigned( 143,8)),
			67 => std_logic_vector(to_unsigned( 43,8)),
			68 => std_logic_vector(to_unsigned( 39,8)),
			69 => std_logic_vector(to_unsigned( 130,8)),
			70 => std_logic_vector(to_unsigned( 75,8)),
			71 => std_logic_vector(to_unsigned( 20,8)),
			72 => std_logic_vector(to_unsigned( 234,8)),
			73 => std_logic_vector(to_unsigned( 113,8)),
			74 => std_logic_vector(to_unsigned( 157,8)),
			75 => std_logic_vector(to_unsigned( 214,8)),
			76 => std_logic_vector(to_unsigned( 183,8)),
			77 => std_logic_vector(to_unsigned( 185,8)),
			78 => std_logic_vector(to_unsigned( 186,8)),
			79 => std_logic_vector(to_unsigned( 123,8)),
			80 => std_logic_vector(to_unsigned( 41,8)),
			81 => std_logic_vector(to_unsigned( 81,8)),
			82 => std_logic_vector(to_unsigned( 180,8)),
			83 => std_logic_vector(to_unsigned( 193,8)),
			84 => std_logic_vector(to_unsigned( 153,8)),
			85 => std_logic_vector(to_unsigned( 68,8)),
			86 => std_logic_vector(to_unsigned( 219,8)),
			87 => std_logic_vector(to_unsigned( 163,8)),
			88 => std_logic_vector(to_unsigned( 252,8)),
			89 => std_logic_vector(to_unsigned( 223,8)),
			90 => std_logic_vector(to_unsigned( 106,8)),
			91 => std_logic_vector(to_unsigned( 184,8)),
			92 => std_logic_vector(to_unsigned( 199,8)),
			93 => std_logic_vector(to_unsigned( 57,8)),
			94 => std_logic_vector(to_unsigned( 111,8)),
			95 => std_logic_vector(to_unsigned( 91,8)),
			96 => std_logic_vector(to_unsigned( 200,8)),
			97 => std_logic_vector(to_unsigned( 155,8)),
			98 => std_logic_vector(to_unsigned( 245,8)),
			99 => std_logic_vector(to_unsigned( 36,8)),
			100 => std_logic_vector(to_unsigned( 141,8)),
			101 => std_logic_vector(to_unsigned( 238,8)),
			102 => std_logic_vector(to_unsigned( 35,8)),
			103 => std_logic_vector(to_unsigned( 74,8)),
			104 => std_logic_vector(to_unsigned( 237,8)),
			105 => std_logic_vector(to_unsigned( 92,8)),
			106 => std_logic_vector(to_unsigned( 207,8)),
			107 => std_logic_vector(to_unsigned( 80,8)),
			108 => std_logic_vector(to_unsigned( 28,8)),
			109 => std_logic_vector(to_unsigned( 10,8)),
			110 => std_logic_vector(to_unsigned( 163,8)),
			111 => std_logic_vector(to_unsigned( 48,8)),
			112 => std_logic_vector(to_unsigned( 127,8)),
			113 => std_logic_vector(to_unsigned( 24,8)),
			114 => std_logic_vector(to_unsigned( 243,8)),
			115 => std_logic_vector(to_unsigned( 185,8)),
			116 => std_logic_vector(to_unsigned( 83,8)),
			117 => std_logic_vector(to_unsigned( 36,8)),
			118 => std_logic_vector(to_unsigned( 241,8)),
			119 => std_logic_vector(to_unsigned( 134,8)),
			120 => std_logic_vector(to_unsigned( 205,8)),
			121 => std_logic_vector(to_unsigned( 87,8)),
			122 => std_logic_vector(to_unsigned( 45,8)),
			123 => std_logic_vector(to_unsigned( 184,8)),
			124 => std_logic_vector(to_unsigned( 52,8)),
			125 => std_logic_vector(to_unsigned( 126,8)),
			126 => std_logic_vector(to_unsigned( 155,8)),
			127 => std_logic_vector(to_unsigned( 41,8)),
			128 => std_logic_vector(to_unsigned( 246,8)),
			129 => std_logic_vector(to_unsigned( 213,8)),
			130 => std_logic_vector(to_unsigned( 123,8)),
			131 => std_logic_vector(to_unsigned( 99,8)),
			132 => std_logic_vector(to_unsigned( 181,8)),
			133 => std_logic_vector(to_unsigned( 215,8)),
			134 => std_logic_vector(to_unsigned( 4,8)),
			135 => std_logic_vector(to_unsigned( 36,8)),
			136 => std_logic_vector(to_unsigned( 169,8)),
			137 => std_logic_vector(to_unsigned( 155,8)),
			138 => std_logic_vector(to_unsigned( 208,8)),
			139 => std_logic_vector(to_unsigned( 128,8)),
			140 => std_logic_vector(to_unsigned( 89,8)),
			141 => std_logic_vector(to_unsigned( 3,8)),
			142 => std_logic_vector(to_unsigned( 151,8)),
			143 => std_logic_vector(to_unsigned( 247,8)),
			144 => std_logic_vector(to_unsigned( 228,8)),
			145 => std_logic_vector(to_unsigned( 17,8)),
			146 => std_logic_vector(to_unsigned( 43,8)),
			147 => std_logic_vector(to_unsigned( 145,8)),
			148 => std_logic_vector(to_unsigned( 35,8)),
			149 => std_logic_vector(to_unsigned( 231,8)),
			150 => std_logic_vector(to_unsigned( 133,8)),
			151 => std_logic_vector(to_unsigned( 191,8)),
			152 => std_logic_vector(to_unsigned( 66,8)),
			153 => std_logic_vector(to_unsigned( 149,8)),
			154 => std_logic_vector(to_unsigned( 77,8)),
			155 => std_logic_vector(to_unsigned( 41,8)),
			156 => std_logic_vector(to_unsigned( 123,8)),
			157 => std_logic_vector(to_unsigned( 97,8)),
			158 => std_logic_vector(to_unsigned( 248,8)),
			159 => std_logic_vector(to_unsigned( 119,8)),
			160 => std_logic_vector(to_unsigned( 58,8)),
			161 => std_logic_vector(to_unsigned( 136,8)),
			162 => std_logic_vector(to_unsigned( 91,8)),
			163 => std_logic_vector(to_unsigned( 40,8)),
			164 => std_logic_vector(to_unsigned( 70,8)),
			165 => std_logic_vector(to_unsigned( 139,8)),
			166 => std_logic_vector(to_unsigned( 10,8)),
			167 => std_logic_vector(to_unsigned( 234,8)),
			168 => std_logic_vector(to_unsigned( 224,8)),
			169 => std_logic_vector(to_unsigned( 194,8)),
			170 => std_logic_vector(to_unsigned( 75,8)),
			171 => std_logic_vector(to_unsigned( 0,8)),
			172 => std_logic_vector(to_unsigned( 226,8)),
			173 => std_logic_vector(to_unsigned( 66,8)),
			174 => std_logic_vector(to_unsigned( 253,8)),
			175 => std_logic_vector(to_unsigned( 87,8)),
			176 => std_logic_vector(to_unsigned( 78,8)),
			177 => std_logic_vector(to_unsigned( 121,8)),
			178 => std_logic_vector(to_unsigned( 200,8)),
			179 => std_logic_vector(to_unsigned( 41,8)),
			180 => std_logic_vector(to_unsigned( 216,8)),
			181 => std_logic_vector(to_unsigned( 227,8)),
			182 => std_logic_vector(to_unsigned( 171,8)),
			183 => std_logic_vector(to_unsigned( 153,8)),
			184 => std_logic_vector(to_unsigned( 158,8)),
			185 => std_logic_vector(to_unsigned( 107,8)),
			186 => std_logic_vector(to_unsigned( 11,8)),
			187 => std_logic_vector(to_unsigned( 108,8)),
			188 => std_logic_vector(to_unsigned( 217,8)),
			189 => std_logic_vector(to_unsigned( 118,8)),
			190 => std_logic_vector(to_unsigned( 104,8)),
			191 => std_logic_vector(to_unsigned( 212,8)),
			192 => std_logic_vector(to_unsigned( 0,8)),
			193 => std_logic_vector(to_unsigned( 80,8)),
			194 => std_logic_vector(to_unsigned( 159,8)),
			195 => std_logic_vector(to_unsigned( 134,8)),
			196 => std_logic_vector(to_unsigned( 192,8)),
			197 => std_logic_vector(to_unsigned( 55,8)),
			198 => std_logic_vector(to_unsigned( 234,8)),
			199 => std_logic_vector(to_unsigned( 50,8)),
			200 => std_logic_vector(to_unsigned( 124,8)),
			201 => std_logic_vector(to_unsigned( 153,8)),
			202 => std_logic_vector(to_unsigned( 226,8)),
			203 => std_logic_vector(to_unsigned( 2,8)),
			204 => std_logic_vector(to_unsigned( 92,8)),
			205 => std_logic_vector(to_unsigned( 88,8)),
			206 => std_logic_vector(to_unsigned( 135,8)),
			207 => std_logic_vector(to_unsigned( 182,8)),
			208 => std_logic_vector(to_unsigned( 92,8)),
			209 => std_logic_vector(to_unsigned( 205,8)),
			210 => std_logic_vector(to_unsigned( 92,8)),
			211 => std_logic_vector(to_unsigned( 42,8)),
			212 => std_logic_vector(to_unsigned( 29,8)),
			213 => std_logic_vector(to_unsigned( 50,8)),
			214 => std_logic_vector(to_unsigned( 188,8)),
			215 => std_logic_vector(to_unsigned( 100,8)),
			216 => std_logic_vector(to_unsigned( 3,8)),
			217 => std_logic_vector(to_unsigned( 47,8)),
			218 => std_logic_vector(to_unsigned( 111,8)),
			219 => std_logic_vector(to_unsigned( 108,8)),
			220 => std_logic_vector(to_unsigned( 72,8)),
			221 => std_logic_vector(to_unsigned( 79,8)),
			222 => std_logic_vector(to_unsigned( 128,8)),
			223 => std_logic_vector(to_unsigned( 11,8)),
			224 => std_logic_vector(to_unsigned( 155,8)),
			225 => std_logic_vector(to_unsigned( 237,8)),
			226 => std_logic_vector(to_unsigned( 165,8)),
			227 => std_logic_vector(to_unsigned( 251,8)),
			228 => std_logic_vector(to_unsigned( 230,8)),
			229 => std_logic_vector(to_unsigned( 136,8)),
			230 => std_logic_vector(to_unsigned( 73,8)),
			231 => std_logic_vector(to_unsigned( 41,8)),
			232 => std_logic_vector(to_unsigned( 190,8)),
			233 => std_logic_vector(to_unsigned( 64,8)),
			234 => std_logic_vector(to_unsigned( 205,8)),
			235 => std_logic_vector(to_unsigned( 165,8)),
			236 => std_logic_vector(to_unsigned( 103,8)),
			237 => std_logic_vector(to_unsigned( 133,8)),
			238 => std_logic_vector(to_unsigned( 204,8)),
			239 => std_logic_vector(to_unsigned( 177,8)),
			240 => std_logic_vector(to_unsigned( 138,8)),
			241 => std_logic_vector(to_unsigned( 17,8)),
			242 => std_logic_vector(to_unsigned( 255,8)),
			243 => std_logic_vector(to_unsigned( 107,8)),
			244 => std_logic_vector(to_unsigned( 250,8)),
			245 => std_logic_vector(to_unsigned( 135,8)),
			246 => std_logic_vector(to_unsigned( 26,8)),
			247 => std_logic_vector(to_unsigned( 154,8)),
			248 => std_logic_vector(to_unsigned( 226,8)),
			249 => std_logic_vector(to_unsigned( 74,8)),
			250 => std_logic_vector(to_unsigned( 5,8)),
			251 => std_logic_vector(to_unsigned( 21,8)),
			252 => std_logic_vector(to_unsigned( 153,8)),
			253 => std_logic_vector(to_unsigned( 121,8)),
			254 => std_logic_vector(to_unsigned( 210,8)),
			255 => std_logic_vector(to_unsigned( 234,8)),
			256 => std_logic_vector(to_unsigned( 235,8)),
			257 => std_logic_vector(to_unsigned( 81,8)),
			258 => std_logic_vector(to_unsigned( 158,8)),
			259 => std_logic_vector(to_unsigned( 37,8)),
			260 => std_logic_vector(to_unsigned( 157,8)),
			261 => std_logic_vector(to_unsigned( 128,8)),
			262 => std_logic_vector(to_unsigned( 244,8)),
			263 => std_logic_vector(to_unsigned( 206,8)),
			264 => std_logic_vector(to_unsigned( 210,8)),
			265 => std_logic_vector(to_unsigned( 7,8)),
			266 => std_logic_vector(to_unsigned( 174,8)),
			267 => std_logic_vector(to_unsigned( 230,8)),
			268 => std_logic_vector(to_unsigned( 95,8)),
			269 => std_logic_vector(to_unsigned( 213,8)),
			270 => std_logic_vector(to_unsigned( 174,8)),
			271 => std_logic_vector(to_unsigned( 149,8)),
			272 => std_logic_vector(to_unsigned( 48,8)),
			273 => std_logic_vector(to_unsigned( 125,8)),
			274 => std_logic_vector(to_unsigned( 213,8)),
			275 => std_logic_vector(to_unsigned( 12,8)),
			276 => std_logic_vector(to_unsigned( 138,8)),
			277 => std_logic_vector(to_unsigned( 55,8)),
			278 => std_logic_vector(to_unsigned( 153,8)),
			279 => std_logic_vector(to_unsigned( 168,8)),
			280 => std_logic_vector(to_unsigned( 231,8)),
			281 => std_logic_vector(to_unsigned( 122,8)),
			282 => std_logic_vector(to_unsigned( 160,8)),
			283 => std_logic_vector(to_unsigned( 74,8)),
			284 => std_logic_vector(to_unsigned( 72,8)),
			285 => std_logic_vector(to_unsigned( 96,8)),
			286 => std_logic_vector(to_unsigned( 214,8)),
			287 => std_logic_vector(to_unsigned( 19,8)),
			288 => std_logic_vector(to_unsigned( 82,8)),
			289 => std_logic_vector(to_unsigned( 134,8)),
			290 => std_logic_vector(to_unsigned( 249,8)),
			291 => std_logic_vector(to_unsigned( 243,8)),
			292 => std_logic_vector(to_unsigned( 224,8)),
			293 => std_logic_vector(to_unsigned( 105,8)),
			294 => std_logic_vector(to_unsigned( 149,8)),
			295 => std_logic_vector(to_unsigned( 184,8)),
			296 => std_logic_vector(to_unsigned( 54,8)),
			297 => std_logic_vector(to_unsigned( 203,8)),
			298 => std_logic_vector(to_unsigned( 122,8)),
			299 => std_logic_vector(to_unsigned( 60,8)),
			300 => std_logic_vector(to_unsigned( 70,8)),
			301 => std_logic_vector(to_unsigned( 138,8)),
			302 => std_logic_vector(to_unsigned( 196,8)),
			303 => std_logic_vector(to_unsigned( 70,8)),
			304 => std_logic_vector(to_unsigned( 203,8)),
			305 => std_logic_vector(to_unsigned( 202,8)),
			306 => std_logic_vector(to_unsigned( 129,8)),
			307 => std_logic_vector(to_unsigned( 153,8)),
			308 => std_logic_vector(to_unsigned( 119,8)),
			309 => std_logic_vector(to_unsigned( 98,8)),
			310 => std_logic_vector(to_unsigned( 57,8)),
			311 => std_logic_vector(to_unsigned( 176,8)),
			312 => std_logic_vector(to_unsigned( 47,8)),
			313 => std_logic_vector(to_unsigned( 224,8)),
			314 => std_logic_vector(to_unsigned( 7,8)),
			315 => std_logic_vector(to_unsigned( 121,8)),
			316 => std_logic_vector(to_unsigned( 38,8)),
			317 => std_logic_vector(to_unsigned( 154,8)),
			318 => std_logic_vector(to_unsigned( 64,8)),
			319 => std_logic_vector(to_unsigned( 209,8)),
			320 => std_logic_vector(to_unsigned( 56,8)),
			321 => std_logic_vector(to_unsigned( 131,8)),
			322 => std_logic_vector(to_unsigned( 221,8)),
			323 => std_logic_vector(to_unsigned( 68,8)),
			324 => std_logic_vector(to_unsigned( 87,8)),
			325 => std_logic_vector(to_unsigned( 97,8)),
			326 => std_logic_vector(to_unsigned( 6,8)),
			327 => std_logic_vector(to_unsigned( 162,8)),
			328 => std_logic_vector(to_unsigned( 233,8)),
			329 => std_logic_vector(to_unsigned( 182,8)),
			330 => std_logic_vector(to_unsigned( 130,8)),
			331 => std_logic_vector(to_unsigned( 193,8)),
			332 => std_logic_vector(to_unsigned( 248,8)),
			333 => std_logic_vector(to_unsigned( 142,8)),
			334 => std_logic_vector(to_unsigned( 171,8)),
			335 => std_logic_vector(to_unsigned( 232,8)),
			336 => std_logic_vector(to_unsigned( 69,8)),
			337 => std_logic_vector(to_unsigned( 0,8)),
			338 => std_logic_vector(to_unsigned( 188,8)),
			339 => std_logic_vector(to_unsigned( 225,8)),
			340 => std_logic_vector(to_unsigned( 35,8)),
			341 => std_logic_vector(to_unsigned( 144,8)),
			342 => std_logic_vector(to_unsigned( 152,8)),
			343 => std_logic_vector(to_unsigned( 251,8)),
			344 => std_logic_vector(to_unsigned( 102,8)),
			345 => std_logic_vector(to_unsigned( 83,8)),
			346 => std_logic_vector(to_unsigned( 111,8)),
			347 => std_logic_vector(to_unsigned( 18,8)),
			348 => std_logic_vector(to_unsigned( 201,8)),
			349 => std_logic_vector(to_unsigned( 224,8)),
			350 => std_logic_vector(to_unsigned( 5,8)),
			351 => std_logic_vector(to_unsigned( 215,8)),
			352 => std_logic_vector(to_unsigned( 93,8)),
			353 => std_logic_vector(to_unsigned( 233,8)),
			354 => std_logic_vector(to_unsigned( 199,8)),
			355 => std_logic_vector(to_unsigned( 142,8)),
			356 => std_logic_vector(to_unsigned( 36,8)),
			357 => std_logic_vector(to_unsigned( 53,8)),
			358 => std_logic_vector(to_unsigned( 170,8)),
			359 => std_logic_vector(to_unsigned( 25,8)),
			360 => std_logic_vector(to_unsigned( 170,8)),
			361 => std_logic_vector(to_unsigned( 3,8)),
			362 => std_logic_vector(to_unsigned( 29,8)),
			363 => std_logic_vector(to_unsigned( 221,8)),
			364 => std_logic_vector(to_unsigned( 65,8)),
			365 => std_logic_vector(to_unsigned( 68,8)),
			366 => std_logic_vector(to_unsigned( 23,8)),
			367 => std_logic_vector(to_unsigned( 245,8)),
			368 => std_logic_vector(to_unsigned( 1,8)),
			369 => std_logic_vector(to_unsigned( 122,8)),
			370 => std_logic_vector(to_unsigned( 177,8)),
			371 => std_logic_vector(to_unsigned( 154,8)),
			372 => std_logic_vector(to_unsigned( 127,8)),
			373 => std_logic_vector(to_unsigned( 225,8)),
			374 => std_logic_vector(to_unsigned( 134,8)),
			375 => std_logic_vector(to_unsigned( 6,8)),
			376 => std_logic_vector(to_unsigned( 209,8)),
			377 => std_logic_vector(to_unsigned( 108,8)),
			378 => std_logic_vector(to_unsigned( 209,8)),
			379 => std_logic_vector(to_unsigned( 119,8)),
			380 => std_logic_vector(to_unsigned( 245,8)),
			381 => std_logic_vector(to_unsigned( 65,8)),
			382 => std_logic_vector(to_unsigned( 166,8)),
			383 => std_logic_vector(to_unsigned( 137,8)),
			384 => std_logic_vector(to_unsigned( 229,8)),
			385 => std_logic_vector(to_unsigned( 194,8)),
			386 => std_logic_vector(to_unsigned( 134,8)),
			387 => std_logic_vector(to_unsigned( 233,8)),
			388 => std_logic_vector(to_unsigned( 130,8)),
			389 => std_logic_vector(to_unsigned( 32,8)),
			390 => std_logic_vector(to_unsigned( 13,8)),
			391 => std_logic_vector(to_unsigned( 33,8)),
			392 => std_logic_vector(to_unsigned( 197,8)),
			393 => std_logic_vector(to_unsigned( 124,8)),
			394 => std_logic_vector(to_unsigned( 50,8)),
			395 => std_logic_vector(to_unsigned( 219,8)),
			396 => std_logic_vector(to_unsigned( 54,8)),
			397 => std_logic_vector(to_unsigned( 97,8)),
			398 => std_logic_vector(to_unsigned( 33,8)),
			399 => std_logic_vector(to_unsigned( 237,8)),
			400 => std_logic_vector(to_unsigned( 15,8)),
			401 => std_logic_vector(to_unsigned( 112,8)),
			402 => std_logic_vector(to_unsigned( 49,8)),
			403 => std_logic_vector(to_unsigned( 253,8)),
			404 => std_logic_vector(to_unsigned( 229,8)),
			405 => std_logic_vector(to_unsigned( 119,8)),
			406 => std_logic_vector(to_unsigned( 44,8)),
			407 => std_logic_vector(to_unsigned( 29,8)),
			408 => std_logic_vector(to_unsigned( 150,8)),
			409 => std_logic_vector(to_unsigned( 101,8)),
			410 => std_logic_vector(to_unsigned( 18,8)),
			411 => std_logic_vector(to_unsigned( 107,8)),
			412 => std_logic_vector(to_unsigned( 202,8)),
			413 => std_logic_vector(to_unsigned( 143,8)),
			414 => std_logic_vector(to_unsigned( 70,8)),
			415 => std_logic_vector(to_unsigned( 244,8)),
			416 => std_logic_vector(to_unsigned( 137,8)),
			417 => std_logic_vector(to_unsigned( 124,8)),
			418 => std_logic_vector(to_unsigned( 188,8)),
			419 => std_logic_vector(to_unsigned( 187,8)),
			420 => std_logic_vector(to_unsigned( 189,8)),
			421 => std_logic_vector(to_unsigned( 130,8)),
			422 => std_logic_vector(to_unsigned( 207,8)),
			423 => std_logic_vector(to_unsigned( 230,8)),
			424 => std_logic_vector(to_unsigned( 254,8)),
			425 => std_logic_vector(to_unsigned( 102,8)),
			426 => std_logic_vector(to_unsigned( 223,8)),
			427 => std_logic_vector(to_unsigned( 44,8)),
			428 => std_logic_vector(to_unsigned( 191,8)),
			429 => std_logic_vector(to_unsigned( 221,8)),
			430 => std_logic_vector(to_unsigned( 218,8)),
			431 => std_logic_vector(to_unsigned( 155,8)),
			432 => std_logic_vector(to_unsigned( 229,8)),
			433 => std_logic_vector(to_unsigned( 93,8)),
			434 => std_logic_vector(to_unsigned( 176,8)),
			435 => std_logic_vector(to_unsigned( 12,8)),
			436 => std_logic_vector(to_unsigned( 111,8)),
			437 => std_logic_vector(to_unsigned( 205,8)),
			438 => std_logic_vector(to_unsigned( 51,8)),
			439 => std_logic_vector(to_unsigned( 217,8)),
			440 => std_logic_vector(to_unsigned( 21,8)),
			441 => std_logic_vector(to_unsigned( 249,8)),
			442 => std_logic_vector(to_unsigned( 202,8)),
			443 => std_logic_vector(to_unsigned( 182,8)),
			444 => std_logic_vector(to_unsigned( 16,8)),
			445 => std_logic_vector(to_unsigned( 38,8)),
			446 => std_logic_vector(to_unsigned( 174,8)),
			447 => std_logic_vector(to_unsigned( 219,8)),
			448 => std_logic_vector(to_unsigned( 61,8)),
			449 => std_logic_vector(to_unsigned( 7,8)),
			450 => std_logic_vector(to_unsigned( 242,8)),
			451 => std_logic_vector(to_unsigned( 167,8)),
			452 => std_logic_vector(to_unsigned( 69,8)),
			453 => std_logic_vector(to_unsigned( 37,8)),
			454 => std_logic_vector(to_unsigned( 221,8)),
			455 => std_logic_vector(to_unsigned( 185,8)),
			456 => std_logic_vector(to_unsigned( 187,8)),
			457 => std_logic_vector(to_unsigned( 86,8)),
			458 => std_logic_vector(to_unsigned( 96,8)),
			459 => std_logic_vector(to_unsigned( 16,8)),
			460 => std_logic_vector(to_unsigned( 174,8)),
			461 => std_logic_vector(to_unsigned( 31,8)),
			462 => std_logic_vector(to_unsigned( 197,8)),
			463 => std_logic_vector(to_unsigned( 177,8)),
			464 => std_logic_vector(to_unsigned( 80,8)),
			465 => std_logic_vector(to_unsigned( 83,8)),
			466 => std_logic_vector(to_unsigned( 200,8)),
			467 => std_logic_vector(to_unsigned( 193,8)),
			468 => std_logic_vector(to_unsigned( 253,8)),
			469 => std_logic_vector(to_unsigned( 28,8)),
			470 => std_logic_vector(to_unsigned( 212,8)),
			471 => std_logic_vector(to_unsigned( 16,8)),
			472 => std_logic_vector(to_unsigned( 47,8)),
			473 => std_logic_vector(to_unsigned( 130,8)),
			474 => std_logic_vector(to_unsigned( 133,8)),
			475 => std_logic_vector(to_unsigned( 24,8)),
			476 => std_logic_vector(to_unsigned( 203,8)),
			477 => std_logic_vector(to_unsigned( 195,8)),
			478 => std_logic_vector(to_unsigned( 69,8)),
			479 => std_logic_vector(to_unsigned( 69,8)),
			480 => std_logic_vector(to_unsigned( 132,8)),
			481 => std_logic_vector(to_unsigned( 73,8)),
			482 => std_logic_vector(to_unsigned( 227,8)),
			483 => std_logic_vector(to_unsigned( 96,8)),
			484 => std_logic_vector(to_unsigned( 86,8)),
			485 => std_logic_vector(to_unsigned( 18,8)),
			486 => std_logic_vector(to_unsigned( 31,8)),
			487 => std_logic_vector(to_unsigned( 98,8)),
			488 => std_logic_vector(to_unsigned( 38,8)),
			489 => std_logic_vector(to_unsigned( 164,8)),
			490 => std_logic_vector(to_unsigned( 9,8)),
			491 => std_logic_vector(to_unsigned( 124,8)),
			492 => std_logic_vector(to_unsigned( 159,8)),
			493 => std_logic_vector(to_unsigned( 101,8)),
			494 => std_logic_vector(to_unsigned( 249,8)),
			495 => std_logic_vector(to_unsigned( 60,8)),
			496 => std_logic_vector(to_unsigned( 175,8)),
			497 => std_logic_vector(to_unsigned( 139,8)),
			498 => std_logic_vector(to_unsigned( 209,8)),
			499 => std_logic_vector(to_unsigned( 110,8)),
			500 => std_logic_vector(to_unsigned( 169,8)),
			501 => std_logic_vector(to_unsigned( 54,8)),
			502 => std_logic_vector(to_unsigned( 117,8)),
			503 => std_logic_vector(to_unsigned( 186,8)),
			504 => std_logic_vector(to_unsigned( 179,8)),
			505 => std_logic_vector(to_unsigned( 87,8)),
			506 => std_logic_vector(to_unsigned( 216,8)),
			507 => std_logic_vector(to_unsigned( 218,8)),
			508 => std_logic_vector(to_unsigned( 216,8)),
			509 => std_logic_vector(to_unsigned( 165,8)),
			510 => std_logic_vector(to_unsigned( 120,8)),
			511 => std_logic_vector(to_unsigned( 253,8)),
			512 => std_logic_vector(to_unsigned( 25,8)),
			513 => std_logic_vector(to_unsigned( 153,8)),
			514 => std_logic_vector(to_unsigned( 231,8)),
			515 => std_logic_vector(to_unsigned( 87,8)),
			516 => std_logic_vector(to_unsigned( 244,8)),
			517 => std_logic_vector(to_unsigned( 218,8)),
			518 => std_logic_vector(to_unsigned( 97,8)),
			519 => std_logic_vector(to_unsigned( 237,8)),
			520 => std_logic_vector(to_unsigned( 40,8)),
			521 => std_logic_vector(to_unsigned( 90,8)),
			522 => std_logic_vector(to_unsigned( 52,8)),
			523 => std_logic_vector(to_unsigned( 100,8)),
			524 => std_logic_vector(to_unsigned( 206,8)),
			525 => std_logic_vector(to_unsigned( 188,8)),
			526 => std_logic_vector(to_unsigned( 227,8)),
			527 => std_logic_vector(to_unsigned( 199,8)),
			528 => std_logic_vector(to_unsigned( 40,8)),
			529 => std_logic_vector(to_unsigned( 6,8)),
			530 => std_logic_vector(to_unsigned( 231,8)),
			531 => std_logic_vector(to_unsigned( 236,8)),
			532 => std_logic_vector(to_unsigned( 25,8)),
			533 => std_logic_vector(to_unsigned( 87,8)),
			534 => std_logic_vector(to_unsigned( 56,8)),
			535 => std_logic_vector(to_unsigned( 81,8)),
			536 => std_logic_vector(to_unsigned( 72,8)),
			537 => std_logic_vector(to_unsigned( 200,8)),
			538 => std_logic_vector(to_unsigned( 108,8)),
			539 => std_logic_vector(to_unsigned( 199,8)),
			540 => std_logic_vector(to_unsigned( 61,8)),
			541 => std_logic_vector(to_unsigned( 123,8)),
			542 => std_logic_vector(to_unsigned( 226,8)),
			543 => std_logic_vector(to_unsigned( 32,8)),
			544 => std_logic_vector(to_unsigned( 38,8)),
			545 => std_logic_vector(to_unsigned( 53,8)),
			546 => std_logic_vector(to_unsigned( 242,8)),
			547 => std_logic_vector(to_unsigned( 164,8)),
			548 => std_logic_vector(to_unsigned( 62,8)),
			549 => std_logic_vector(to_unsigned( 231,8)),
			550 => std_logic_vector(to_unsigned( 194,8)),
			551 => std_logic_vector(to_unsigned( 87,8)),
			552 => std_logic_vector(to_unsigned( 246,8)),
			553 => std_logic_vector(to_unsigned( 115,8)),
			554 => std_logic_vector(to_unsigned( 133,8)),
			555 => std_logic_vector(to_unsigned( 39,8)),
			556 => std_logic_vector(to_unsigned( 242,8)),
			557 => std_logic_vector(to_unsigned( 27,8)),
			558 => std_logic_vector(to_unsigned( 18,8)),
			559 => std_logic_vector(to_unsigned( 91,8)),
			560 => std_logic_vector(to_unsigned( 36,8)),
			561 => std_logic_vector(to_unsigned( 115,8)),
			562 => std_logic_vector(to_unsigned( 186,8)),
			563 => std_logic_vector(to_unsigned( 156,8)),
			564 => std_logic_vector(to_unsigned( 107,8)),
			565 => std_logic_vector(to_unsigned( 3,8)),
			566 => std_logic_vector(to_unsigned( 200,8)),
			567 => std_logic_vector(to_unsigned( 227,8)),
			568 => std_logic_vector(to_unsigned( 186,8)),
			569 => std_logic_vector(to_unsigned( 35,8)),
			570 => std_logic_vector(to_unsigned( 56,8)),
			571 => std_logic_vector(to_unsigned( 86,8)),
			572 => std_logic_vector(to_unsigned( 18,8)),
			573 => std_logic_vector(to_unsigned( 171,8)),
			574 => std_logic_vector(to_unsigned( 212,8)),
			575 => std_logic_vector(to_unsigned( 142,8)),
			576 => std_logic_vector(to_unsigned( 171,8)),
			577 => std_logic_vector(to_unsigned( 216,8)),
			578 => std_logic_vector(to_unsigned( 70,8)),
			579 => std_logic_vector(to_unsigned( 8,8)),
			580 => std_logic_vector(to_unsigned( 128,8)),
			581 => std_logic_vector(to_unsigned( 67,8)),
			582 => std_logic_vector(to_unsigned( 188,8)),
			583 => std_logic_vector(to_unsigned( 211,8)),
			584 => std_logic_vector(to_unsigned( 250,8)),
			585 => std_logic_vector(to_unsigned( 58,8)),
			586 => std_logic_vector(to_unsigned( 17,8)),
			587 => std_logic_vector(to_unsigned( 192,8)),
			588 => std_logic_vector(to_unsigned( 184,8)),
			589 => std_logic_vector(to_unsigned( 175,8)),
			590 => std_logic_vector(to_unsigned( 197,8)),
			591 => std_logic_vector(to_unsigned( 82,8)),
			592 => std_logic_vector(to_unsigned( 93,8)),
			593 => std_logic_vector(to_unsigned( 33,8)),
			594 => std_logic_vector(to_unsigned( 159,8)),
			595 => std_logic_vector(to_unsigned( 142,8)),
			596 => std_logic_vector(to_unsigned( 100,8)),
			597 => std_logic_vector(to_unsigned( 185,8)),
			598 => std_logic_vector(to_unsigned( 136,8)),
			599 => std_logic_vector(to_unsigned( 162,8)),
			600 => std_logic_vector(to_unsigned( 66,8)),
			601 => std_logic_vector(to_unsigned( 37,8)),
			602 => std_logic_vector(to_unsigned( 157,8)),
			603 => std_logic_vector(to_unsigned( 124,8)),
			604 => std_logic_vector(to_unsigned( 165,8)),
			605 => std_logic_vector(to_unsigned( 104,8)),
			606 => std_logic_vector(to_unsigned( 245,8)),
			607 => std_logic_vector(to_unsigned( 251,8)),
			608 => std_logic_vector(to_unsigned( 126,8)),
			609 => std_logic_vector(to_unsigned( 229,8)),
			610 => std_logic_vector(to_unsigned( 139,8)),
			611 => std_logic_vector(to_unsigned( 78,8)),
			612 => std_logic_vector(to_unsigned( 44,8)),
			613 => std_logic_vector(to_unsigned( 248,8)),
			614 => std_logic_vector(to_unsigned( 185,8)),
			615 => std_logic_vector(to_unsigned( 136,8)),
			616 => std_logic_vector(to_unsigned( 25,8)),
			617 => std_logic_vector(to_unsigned( 32,8)),
			618 => std_logic_vector(to_unsigned( 195,8)),
			619 => std_logic_vector(to_unsigned( 197,8)),
			620 => std_logic_vector(to_unsigned( 124,8)),
			621 => std_logic_vector(to_unsigned( 177,8)),
			622 => std_logic_vector(to_unsigned( 196,8)),
			623 => std_logic_vector(to_unsigned( 191,8)),
			624 => std_logic_vector(to_unsigned( 255,8)),
			625 => std_logic_vector(to_unsigned( 142,8)),
			626 => std_logic_vector(to_unsigned( 155,8)),
			627 => std_logic_vector(to_unsigned( 54,8)),
			628 => std_logic_vector(to_unsigned( 202,8)),
			629 => std_logic_vector(to_unsigned( 30,8)),
			630 => std_logic_vector(to_unsigned( 238,8)),
			631 => std_logic_vector(to_unsigned( 194,8)),
			632 => std_logic_vector(to_unsigned( 222,8)),
			633 => std_logic_vector(to_unsigned( 45,8)),
			634 => std_logic_vector(to_unsigned( 76,8)),
			635 => std_logic_vector(to_unsigned( 197,8)),
			636 => std_logic_vector(to_unsigned( 187,8)),
			637 => std_logic_vector(to_unsigned( 90,8)),
			638 => std_logic_vector(to_unsigned( 119,8)),
			639 => std_logic_vector(to_unsigned( 89,8)),
			640 => std_logic_vector(to_unsigned( 120,8)),
			641 => std_logic_vector(to_unsigned( 112,8)),
			642 => std_logic_vector(to_unsigned( 139,8)),
			643 => std_logic_vector(to_unsigned( 65,8)),
			644 => std_logic_vector(to_unsigned( 35,8)),
			645 => std_logic_vector(to_unsigned( 104,8)),
			646 => std_logic_vector(to_unsigned( 233,8)),
			647 => std_logic_vector(to_unsigned( 35,8)),
			648 => std_logic_vector(to_unsigned( 71,8)),
			649 => std_logic_vector(to_unsigned( 6,8)),
			650 => std_logic_vector(to_unsigned( 48,8)),
			651 => std_logic_vector(to_unsigned( 188,8)),
			652 => std_logic_vector(to_unsigned( 35,8)),
			653 => std_logic_vector(to_unsigned( 209,8)),
			654 => std_logic_vector(to_unsigned( 130,8)),
			655 => std_logic_vector(to_unsigned( 11,8)),
			656 => std_logic_vector(to_unsigned( 33,8)),
			657 => std_logic_vector(to_unsigned( 167,8)),
			658 => std_logic_vector(to_unsigned( 221,8)),
			659 => std_logic_vector(to_unsigned( 202,8)),
			660 => std_logic_vector(to_unsigned( 119,8)),
			661 => std_logic_vector(to_unsigned( 162,8)),
			662 => std_logic_vector(to_unsigned( 139,8)),
			663 => std_logic_vector(to_unsigned( 157,8)),
			664 => std_logic_vector(to_unsigned( 22,8)),
			665 => std_logic_vector(to_unsigned( 82,8)),
			666 => std_logic_vector(to_unsigned( 107,8)),
			667 => std_logic_vector(to_unsigned( 234,8)),
			668 => std_logic_vector(to_unsigned( 155,8)),
			669 => std_logic_vector(to_unsigned( 127,8)),
			670 => std_logic_vector(to_unsigned( 11,8)),
			671 => std_logic_vector(to_unsigned( 189,8)),
			672 => std_logic_vector(to_unsigned( 172,8)),
			673 => std_logic_vector(to_unsigned( 212,8)),
			674 => std_logic_vector(to_unsigned( 106,8)),
			675 => std_logic_vector(to_unsigned( 34,8)),
			676 => std_logic_vector(to_unsigned( 214,8)),
			677 => std_logic_vector(to_unsigned( 110,8)),
			678 => std_logic_vector(to_unsigned( 124,8)),
			679 => std_logic_vector(to_unsigned( 200,8)),
			680 => std_logic_vector(to_unsigned( 6,8)),
			681 => std_logic_vector(to_unsigned( 3,8)),
			682 => std_logic_vector(to_unsigned( 52,8)),
			683 => std_logic_vector(to_unsigned( 246,8)),
			684 => std_logic_vector(to_unsigned( 114,8)),
			685 => std_logic_vector(to_unsigned( 13,8)),
			686 => std_logic_vector(to_unsigned( 211,8)),
			687 => std_logic_vector(to_unsigned( 53,8)),
			688 => std_logic_vector(to_unsigned( 30,8)),
			689 => std_logic_vector(to_unsigned( 24,8)),
			690 => std_logic_vector(to_unsigned( 65,8)),
			691 => std_logic_vector(to_unsigned( 95,8)),
			692 => std_logic_vector(to_unsigned( 132,8)),
			693 => std_logic_vector(to_unsigned( 251,8)),
			694 => std_logic_vector(to_unsigned( 198,8)),
			695 => std_logic_vector(to_unsigned( 193,8)),
			696 => std_logic_vector(to_unsigned( 2,8)),
			697 => std_logic_vector(to_unsigned( 179,8)),
			698 => std_logic_vector(to_unsigned( 203,8)),
			699 => std_logic_vector(to_unsigned( 85,8)),
			700 => std_logic_vector(to_unsigned( 79,8)),
			701 => std_logic_vector(to_unsigned( 201,8)),
			702 => std_logic_vector(to_unsigned( 237,8)),
			703 => std_logic_vector(to_unsigned( 106,8)),
			704 => std_logic_vector(to_unsigned( 118,8)),
			705 => std_logic_vector(to_unsigned( 168,8)),
			706 => std_logic_vector(to_unsigned( 6,8)),
			707 => std_logic_vector(to_unsigned( 231,8)),
			708 => std_logic_vector(to_unsigned( 192,8)),
			709 => std_logic_vector(to_unsigned( 24,8)),
			710 => std_logic_vector(to_unsigned( 1,8)),
			711 => std_logic_vector(to_unsigned( 47,8)),
			712 => std_logic_vector(to_unsigned( 112,8)),
			713 => std_logic_vector(to_unsigned( 222,8)),
			714 => std_logic_vector(to_unsigned( 27,8)),
			715 => std_logic_vector(to_unsigned( 150,8)),
			716 => std_logic_vector(to_unsigned( 146,8)),
			717 => std_logic_vector(to_unsigned( 13,8)),
			718 => std_logic_vector(to_unsigned( 176,8)),
			719 => std_logic_vector(to_unsigned( 111,8)),
			720 => std_logic_vector(to_unsigned( 189,8)),
			721 => std_logic_vector(to_unsigned( 223,8)),
			722 => std_logic_vector(to_unsigned( 118,8)),
			723 => std_logic_vector(to_unsigned( 99,8)),
			724 => std_logic_vector(to_unsigned( 234,8)),
			725 => std_logic_vector(to_unsigned( 128,8)),
			726 => std_logic_vector(to_unsigned( 198,8)),
			727 => std_logic_vector(to_unsigned( 98,8)),
			728 => std_logic_vector(to_unsigned( 19,8)),
			729 => std_logic_vector(to_unsigned( 188,8)),
			730 => std_logic_vector(to_unsigned( 60,8)),
			731 => std_logic_vector(to_unsigned( 155,8)),
			732 => std_logic_vector(to_unsigned( 244,8)),
			733 => std_logic_vector(to_unsigned( 205,8)),
			734 => std_logic_vector(to_unsigned( 187,8)),
			735 => std_logic_vector(to_unsigned( 255,8)),
			736 => std_logic_vector(to_unsigned( 68,8)),
			737 => std_logic_vector(to_unsigned( 12,8)),
			738 => std_logic_vector(to_unsigned( 196,8)),
			739 => std_logic_vector(to_unsigned( 243,8)),
			740 => std_logic_vector(to_unsigned( 183,8)),
			741 => std_logic_vector(to_unsigned( 97,8)),
			742 => std_logic_vector(to_unsigned( 121,8)),
			743 => std_logic_vector(to_unsigned( 196,8)),
			744 => std_logic_vector(to_unsigned( 142,8)),
			745 => std_logic_vector(to_unsigned( 227,8)),
			746 => std_logic_vector(to_unsigned( 59,8)),
			747 => std_logic_vector(to_unsigned( 86,8)),
			748 => std_logic_vector(to_unsigned( 241,8)),
			749 => std_logic_vector(to_unsigned( 126,8)),
			750 => std_logic_vector(to_unsigned( 134,8)),
			751 => std_logic_vector(to_unsigned( 21,8)),
			752 => std_logic_vector(to_unsigned( 255,8)),
			753 => std_logic_vector(to_unsigned( 85,8)),
			754 => std_logic_vector(to_unsigned( 179,8)),
			755 => std_logic_vector(to_unsigned( 244,8)),
			756 => std_logic_vector(to_unsigned( 50,8)),
			757 => std_logic_vector(to_unsigned( 55,8)),
			758 => std_logic_vector(to_unsigned( 201,8)),
			759 => std_logic_vector(to_unsigned( 104,8)),
			760 => std_logic_vector(to_unsigned( 80,8)),
			761 => std_logic_vector(to_unsigned( 30,8)),
			762 => std_logic_vector(to_unsigned( 123,8)),
			763 => std_logic_vector(to_unsigned( 10,8)),
			764 => std_logic_vector(to_unsigned( 255,8)),
			765 => std_logic_vector(to_unsigned( 54,8)),
			766 => std_logic_vector(to_unsigned( 79,8)),
			767 => std_logic_vector(to_unsigned( 203,8)),
			768 => std_logic_vector(to_unsigned( 89,8)),
			769 => std_logic_vector(to_unsigned( 15,8)),
			770 => std_logic_vector(to_unsigned( 49,8)),
			771 => std_logic_vector(to_unsigned( 135,8)),
			772 => std_logic_vector(to_unsigned( 99,8)),
			773 => std_logic_vector(to_unsigned( 203,8)),
			774 => std_logic_vector(to_unsigned( 16,8)),
			775 => std_logic_vector(to_unsigned( 53,8)),
			776 => std_logic_vector(to_unsigned( 142,8)),
			777 => std_logic_vector(to_unsigned( 111,8)),
			778 => std_logic_vector(to_unsigned( 141,8)),
			779 => std_logic_vector(to_unsigned( 243,8)),
			780 => std_logic_vector(to_unsigned( 138,8)),
			781 => std_logic_vector(to_unsigned( 93,8)),
			782 => std_logic_vector(to_unsigned( 120,8)),
			783 => std_logic_vector(to_unsigned( 156,8)),
			784 => std_logic_vector(to_unsigned( 63,8)),
			785 => std_logic_vector(to_unsigned( 58,8)),
			786 => std_logic_vector(to_unsigned( 117,8)),
			787 => std_logic_vector(to_unsigned( 24,8)),
			788 => std_logic_vector(to_unsigned( 48,8)),
			789 => std_logic_vector(to_unsigned( 161,8)),
			790 => std_logic_vector(to_unsigned( 142,8)),
			791 => std_logic_vector(to_unsigned( 11,8)),
			792 => std_logic_vector(to_unsigned( 247,8)),
			793 => std_logic_vector(to_unsigned( 55,8)),
			794 => std_logic_vector(to_unsigned( 14,8)),
			795 => std_logic_vector(to_unsigned( 161,8)),
			796 => std_logic_vector(to_unsigned( 168,8)),
			797 => std_logic_vector(to_unsigned( 72,8)),
			798 => std_logic_vector(to_unsigned( 140,8)),
			799 => std_logic_vector(to_unsigned( 163,8)),
			800 => std_logic_vector(to_unsigned( 233,8)),
			801 => std_logic_vector(to_unsigned( 79,8)),
			802 => std_logic_vector(to_unsigned( 255,8)),
			803 => std_logic_vector(to_unsigned( 26,8)),
			804 => std_logic_vector(to_unsigned( 115,8)),
			805 => std_logic_vector(to_unsigned( 221,8)),
			806 => std_logic_vector(to_unsigned( 159,8)),
			807 => std_logic_vector(to_unsigned( 54,8)),
			808 => std_logic_vector(to_unsigned( 127,8)),
			809 => std_logic_vector(to_unsigned( 59,8)),
			810 => std_logic_vector(to_unsigned( 29,8)),
			811 => std_logic_vector(to_unsigned( 42,8)),
			812 => std_logic_vector(to_unsigned( 241,8)),
			813 => std_logic_vector(to_unsigned( 72,8)),
			814 => std_logic_vector(to_unsigned( 3,8)),
			815 => std_logic_vector(to_unsigned( 44,8)),
			816 => std_logic_vector(to_unsigned( 7,8)),
			817 => std_logic_vector(to_unsigned( 207,8)),
			818 => std_logic_vector(to_unsigned( 134,8)),
			819 => std_logic_vector(to_unsigned( 25,8)),
			820 => std_logic_vector(to_unsigned( 215,8)),
			821 => std_logic_vector(to_unsigned( 106,8)),
			822 => std_logic_vector(to_unsigned( 124,8)),
			823 => std_logic_vector(to_unsigned( 30,8)),
			824 => std_logic_vector(to_unsigned( 146,8)),
			825 => std_logic_vector(to_unsigned( 221,8)),
			826 => std_logic_vector(to_unsigned( 120,8)),
			827 => std_logic_vector(to_unsigned( 4,8)),
			828 => std_logic_vector(to_unsigned( 76,8)),
			829 => std_logic_vector(to_unsigned( 89,8)),
			830 => std_logic_vector(to_unsigned( 88,8)),
			831 => std_logic_vector(to_unsigned( 1,8)),
			832 => std_logic_vector(to_unsigned( 78,8)),
			833 => std_logic_vector(to_unsigned( 182,8)),
			834 => std_logic_vector(to_unsigned( 144,8)),
			835 => std_logic_vector(to_unsigned( 36,8)),
			836 => std_logic_vector(to_unsigned( 96,8)),
			837 => std_logic_vector(to_unsigned( 143,8)),
			838 => std_logic_vector(to_unsigned( 97,8)),
			839 => std_logic_vector(to_unsigned( 218,8)),
			840 => std_logic_vector(to_unsigned( 39,8)),
			841 => std_logic_vector(to_unsigned( 240,8)),
			842 => std_logic_vector(to_unsigned( 66,8)),
			843 => std_logic_vector(to_unsigned( 59,8)),
			844 => std_logic_vector(to_unsigned( 43,8)),
			845 => std_logic_vector(to_unsigned( 99,8)),
			846 => std_logic_vector(to_unsigned( 131,8)),
			847 => std_logic_vector(to_unsigned( 120,8)),
			848 => std_logic_vector(to_unsigned( 182,8)),
			849 => std_logic_vector(to_unsigned( 109,8)),
			850 => std_logic_vector(to_unsigned( 43,8)),
			851 => std_logic_vector(to_unsigned( 17,8)),
			852 => std_logic_vector(to_unsigned( 233,8)),
			853 => std_logic_vector(to_unsigned( 223,8)),
			854 => std_logic_vector(to_unsigned( 11,8)),
			855 => std_logic_vector(to_unsigned( 255,8)),
			856 => std_logic_vector(to_unsigned( 126,8)),
			857 => std_logic_vector(to_unsigned( 216,8)),
			858 => std_logic_vector(to_unsigned( 89,8)),
			859 => std_logic_vector(to_unsigned( 216,8)),
			860 => std_logic_vector(to_unsigned( 67,8)),
			861 => std_logic_vector(to_unsigned( 250,8)),
			862 => std_logic_vector(to_unsigned( 1,8)),
			863 => std_logic_vector(to_unsigned( 5,8)),
			864 => std_logic_vector(to_unsigned( 68,8)),
			865 => std_logic_vector(to_unsigned( 86,8)),
			866 => std_logic_vector(to_unsigned( 211,8)),
			867 => std_logic_vector(to_unsigned( 208,8)),
			868 => std_logic_vector(to_unsigned( 215,8)),
			869 => std_logic_vector(to_unsigned( 249,8)),
			870 => std_logic_vector(to_unsigned( 219,8)),
			871 => std_logic_vector(to_unsigned( 23,8)),
			872 => std_logic_vector(to_unsigned( 126,8)),
			873 => std_logic_vector(to_unsigned( 101,8)),
			874 => std_logic_vector(to_unsigned( 215,8)),
			875 => std_logic_vector(to_unsigned( 105,8)),
			876 => std_logic_vector(to_unsigned( 35,8)),
			877 => std_logic_vector(to_unsigned( 183,8)),
			878 => std_logic_vector(to_unsigned( 64,8)),
			879 => std_logic_vector(to_unsigned( 73,8)),
			880 => std_logic_vector(to_unsigned( 27,8)),
			881 => std_logic_vector(to_unsigned( 34,8)),
			882 => std_logic_vector(to_unsigned( 245,8)),
			883 => std_logic_vector(to_unsigned( 55,8)),
			884 => std_logic_vector(to_unsigned( 114,8)),
			885 => std_logic_vector(to_unsigned( 206,8)),
			886 => std_logic_vector(to_unsigned( 33,8)),
			887 => std_logic_vector(to_unsigned( 147,8)),
			888 => std_logic_vector(to_unsigned( 159,8)),
			889 => std_logic_vector(to_unsigned( 181,8)),
			890 => std_logic_vector(to_unsigned( 99,8)),
			891 => std_logic_vector(to_unsigned( 96,8)),
			892 => std_logic_vector(to_unsigned( 100,8)),
			893 => std_logic_vector(to_unsigned( 123,8)),
			894 => std_logic_vector(to_unsigned( 162,8)),
			895 => std_logic_vector(to_unsigned( 131,8)),
			896 => std_logic_vector(to_unsigned( 91,8)),
			897 => std_logic_vector(to_unsigned( 17,8)),
			898 => std_logic_vector(to_unsigned( 115,8)),
			899 => std_logic_vector(to_unsigned( 66,8)),
			900 => std_logic_vector(to_unsigned( 23,8)),
			901 => std_logic_vector(to_unsigned( 141,8)),
			902 => std_logic_vector(to_unsigned( 122,8)),
			903 => std_logic_vector(to_unsigned( 109,8)),
			904 => std_logic_vector(to_unsigned( 203,8)),
			905 => std_logic_vector(to_unsigned( 35,8)),
			906 => std_logic_vector(to_unsigned( 197,8)),
			907 => std_logic_vector(to_unsigned( 146,8)),
			908 => std_logic_vector(to_unsigned( 14,8)),
			909 => std_logic_vector(to_unsigned( 185,8)),
			910 => std_logic_vector(to_unsigned( 36,8)),
			911 => std_logic_vector(to_unsigned( 254,8)),
			912 => std_logic_vector(to_unsigned( 215,8)),
			913 => std_logic_vector(to_unsigned( 146,8)),
			914 => std_logic_vector(to_unsigned( 208,8)),
			915 => std_logic_vector(to_unsigned( 176,8)),
			916 => std_logic_vector(to_unsigned( 169,8)),
			917 => std_logic_vector(to_unsigned( 192,8)),
			918 => std_logic_vector(to_unsigned( 107,8)),
			919 => std_logic_vector(to_unsigned( 59,8)),
			920 => std_logic_vector(to_unsigned( 239,8)),
			921 => std_logic_vector(to_unsigned( 152,8)),
			922 => std_logic_vector(to_unsigned( 142,8)),
			923 => std_logic_vector(to_unsigned( 56,8)),
			924 => std_logic_vector(to_unsigned( 127,8)),
			925 => std_logic_vector(to_unsigned( 174,8)),
			926 => std_logic_vector(to_unsigned( 188,8)),
			927 => std_logic_vector(to_unsigned( 152,8)),
			928 => std_logic_vector(to_unsigned( 244,8)),
			929 => std_logic_vector(to_unsigned( 219,8)),
			930 => std_logic_vector(to_unsigned( 115,8)),
			931 => std_logic_vector(to_unsigned( 65,8)),
			932 => std_logic_vector(to_unsigned( 169,8)),
			933 => std_logic_vector(to_unsigned( 75,8)),
			934 => std_logic_vector(to_unsigned( 186,8)),
			935 => std_logic_vector(to_unsigned( 122,8)),
			936 => std_logic_vector(to_unsigned( 62,8)),
			937 => std_logic_vector(to_unsigned( 205,8)),
			938 => std_logic_vector(to_unsigned( 157,8)),
			939 => std_logic_vector(to_unsigned( 113,8)),
			940 => std_logic_vector(to_unsigned( 70,8)),
			941 => std_logic_vector(to_unsigned( 11,8)),
			942 => std_logic_vector(to_unsigned( 183,8)),
			943 => std_logic_vector(to_unsigned( 247,8)),
			944 => std_logic_vector(to_unsigned( 234,8)),
			945 => std_logic_vector(to_unsigned( 109,8)),
			946 => std_logic_vector(to_unsigned( 175,8)),
			947 => std_logic_vector(to_unsigned( 185,8)),
			948 => std_logic_vector(to_unsigned( 250,8)),
			949 => std_logic_vector(to_unsigned( 172,8)),
			950 => std_logic_vector(to_unsigned( 189,8)),
			951 => std_logic_vector(to_unsigned( 139,8)),
			952 => std_logic_vector(to_unsigned( 3,8)),
			953 => std_logic_vector(to_unsigned( 140,8)),
			954 => std_logic_vector(to_unsigned( 202,8)),
			955 => std_logic_vector(to_unsigned( 142,8)),
			956 => std_logic_vector(to_unsigned( 99,8)),
			957 => std_logic_vector(to_unsigned( 52,8)),
			958 => std_logic_vector(to_unsigned( 207,8)),
			959 => std_logic_vector(to_unsigned( 225,8)),
			960 => std_logic_vector(to_unsigned( 89,8)),
			961 => std_logic_vector(to_unsigned( 246,8)),
			962 => std_logic_vector(to_unsigned( 115,8)),
			963 => std_logic_vector(to_unsigned( 73,8)),
			964 => std_logic_vector(to_unsigned( 91,8)),
			965 => std_logic_vector(to_unsigned( 139,8)),
			966 => std_logic_vector(to_unsigned( 176,8)),
			967 => std_logic_vector(to_unsigned( 121,8)),
			968 => std_logic_vector(to_unsigned( 195,8)),
			969 => std_logic_vector(to_unsigned( 72,8)),
			970 => std_logic_vector(to_unsigned( 89,8)),
			971 => std_logic_vector(to_unsigned( 83,8)),
			972 => std_logic_vector(to_unsigned( 145,8)),
			973 => std_logic_vector(to_unsigned( 121,8)),
			974 => std_logic_vector(to_unsigned( 30,8)),
			975 => std_logic_vector(to_unsigned( 145,8)),
			976 => std_logic_vector(to_unsigned( 195,8)),
			977 => std_logic_vector(to_unsigned( 155,8)),
			978 => std_logic_vector(to_unsigned( 177,8)),
			979 => std_logic_vector(to_unsigned( 185,8)),
			980 => std_logic_vector(to_unsigned( 79,8)),
			981 => std_logic_vector(to_unsigned( 7,8)),
			982 => std_logic_vector(to_unsigned( 114,8)),
			983 => std_logic_vector(to_unsigned( 225,8)),
			984 => std_logic_vector(to_unsigned( 245,8)),
			985 => std_logic_vector(to_unsigned( 118,8)),
			986 => std_logic_vector(to_unsigned( 222,8)),
			987 => std_logic_vector(to_unsigned( 211,8)),
			988 => std_logic_vector(to_unsigned( 195,8)),
			989 => std_logic_vector(to_unsigned( 96,8)),
			990 => std_logic_vector(to_unsigned( 129,8)),
			991 => std_logic_vector(to_unsigned( 188,8)),
			992 => std_logic_vector(to_unsigned( 118,8)),
			993 => std_logic_vector(to_unsigned( 253,8)),
			994 => std_logic_vector(to_unsigned( 97,8)),
			995 => std_logic_vector(to_unsigned( 202,8)),
			996 => std_logic_vector(to_unsigned( 155,8)),
			997 => std_logic_vector(to_unsigned( 56,8)),
			998 => std_logic_vector(to_unsigned( 201,8)),
			999 => std_logic_vector(to_unsigned( 50,8)),
			1000 => std_logic_vector(to_unsigned( 36,8)),
			1001 => std_logic_vector(to_unsigned( 216,8)),
			1002 => std_logic_vector(to_unsigned( 37,8)),
			1003 => std_logic_vector(to_unsigned( 219,8)),
			1004 => std_logic_vector(to_unsigned( 175,8)),
			1005 => std_logic_vector(to_unsigned( 94,8)),
			1006 => std_logic_vector(to_unsigned( 242,8)),
			1007 => std_logic_vector(to_unsigned( 29,8)),
			1008 => std_logic_vector(to_unsigned( 150,8)),
			1009 => std_logic_vector(to_unsigned( 232,8)),
			1010 => std_logic_vector(to_unsigned( 226,8)),
			1011 => std_logic_vector(to_unsigned( 195,8)),
			1012 => std_logic_vector(to_unsigned( 87,8)),
			1013 => std_logic_vector(to_unsigned( 122,8)),
			1014 => std_logic_vector(to_unsigned( 210,8)),
			1015 => std_logic_vector(to_unsigned( 239,8)),
			1016 => std_logic_vector(to_unsigned( 21,8)),
			1017 => std_logic_vector(to_unsigned( 220,8)),
			1018 => std_logic_vector(to_unsigned( 27,8)),
			1019 => std_logic_vector(to_unsigned( 228,8)),
			1020 => std_logic_vector(to_unsigned( 59,8)),
			1021 => std_logic_vector(to_unsigned( 162,8)),
			1022 => std_logic_vector(to_unsigned( 92,8)),
			1023 => std_logic_vector(to_unsigned( 215,8)),
			1024 => std_logic_vector(to_unsigned( 254,8)),
			1025 => std_logic_vector(to_unsigned( 59,8)),
			1026 => std_logic_vector(to_unsigned( 62,8)),
			1027 => std_logic_vector(to_unsigned( 78,8)),
			1028 => std_logic_vector(to_unsigned( 194,8)),
			1029 => std_logic_vector(to_unsigned( 189,8)),
			1030 => std_logic_vector(to_unsigned( 53,8)),
			1031 => std_logic_vector(to_unsigned( 27,8)),
			1032 => std_logic_vector(to_unsigned( 143,8)),
			1033 => std_logic_vector(to_unsigned( 228,8)),
			1034 => std_logic_vector(to_unsigned( 169,8)),
			1035 => std_logic_vector(to_unsigned( 164,8)),
			1036 => std_logic_vector(to_unsigned( 43,8)),
			1037 => std_logic_vector(to_unsigned( 100,8)),
			1038 => std_logic_vector(to_unsigned( 248,8)),
			1039 => std_logic_vector(to_unsigned( 9,8)),
			1040 => std_logic_vector(to_unsigned( 159,8)),
			1041 => std_logic_vector(to_unsigned( 69,8)),
			1042 => std_logic_vector(to_unsigned( 37,8)),
			1043 => std_logic_vector(to_unsigned( 44,8)),
			1044 => std_logic_vector(to_unsigned( 66,8)),
			1045 => std_logic_vector(to_unsigned( 92,8)),
			1046 => std_logic_vector(to_unsigned( 73,8)),
			1047 => std_logic_vector(to_unsigned( 89,8)),
			1048 => std_logic_vector(to_unsigned( 230,8)),
			1049 => std_logic_vector(to_unsigned( 112,8)),
			1050 => std_logic_vector(to_unsigned( 181,8)),
			1051 => std_logic_vector(to_unsigned( 35,8)),
			1052 => std_logic_vector(to_unsigned( 95,8)),
			1053 => std_logic_vector(to_unsigned( 255,8)),
			1054 => std_logic_vector(to_unsigned( 234,8)),
			1055 => std_logic_vector(to_unsigned( 174,8)),
			1056 => std_logic_vector(to_unsigned( 6,8)),
			1057 => std_logic_vector(to_unsigned( 59,8)),
			1058 => std_logic_vector(to_unsigned( 73,8)),
			1059 => std_logic_vector(to_unsigned( 108,8)),
			1060 => std_logic_vector(to_unsigned( 228,8)),
			1061 => std_logic_vector(to_unsigned( 57,8)),
			1062 => std_logic_vector(to_unsigned( 166,8)),
			1063 => std_logic_vector(to_unsigned( 144,8)),
			1064 => std_logic_vector(to_unsigned( 84,8)),
			1065 => std_logic_vector(to_unsigned( 94,8)),
			1066 => std_logic_vector(to_unsigned( 31,8)),
			1067 => std_logic_vector(to_unsigned( 123,8)),
			1068 => std_logic_vector(to_unsigned( 115,8)),
			1069 => std_logic_vector(to_unsigned( 190,8)),
			1070 => std_logic_vector(to_unsigned( 242,8)),
			1071 => std_logic_vector(to_unsigned( 187,8)),
			1072 => std_logic_vector(to_unsigned( 161,8)),
			1073 => std_logic_vector(to_unsigned( 231,8)),
			1074 => std_logic_vector(to_unsigned( 220,8)),
			1075 => std_logic_vector(to_unsigned( 250,8)),
			1076 => std_logic_vector(to_unsigned( 97,8)),
			1077 => std_logic_vector(to_unsigned( 215,8)),
			1078 => std_logic_vector(to_unsigned( 177,8)),
			1079 => std_logic_vector(to_unsigned( 69,8)),
			1080 => std_logic_vector(to_unsigned( 52,8)),
			1081 => std_logic_vector(to_unsigned( 137,8)),
			1082 => std_logic_vector(to_unsigned( 117,8)),
			1083 => std_logic_vector(to_unsigned( 143,8)),
			1084 => std_logic_vector(to_unsigned( 55,8)),
			1085 => std_logic_vector(to_unsigned( 36,8)),
			1086 => std_logic_vector(to_unsigned( 118,8)),
			1087 => std_logic_vector(to_unsigned( 80,8)),
			1088 => std_logic_vector(to_unsigned( 213,8)),
			1089 => std_logic_vector(to_unsigned( 167,8)),
			1090 => std_logic_vector(to_unsigned( 206,8)),
			1091 => std_logic_vector(to_unsigned( 17,8)),
			1092 => std_logic_vector(to_unsigned( 109,8)),
			1093 => std_logic_vector(to_unsigned( 6,8)),
			1094 => std_logic_vector(to_unsigned( 162,8)),
			1095 => std_logic_vector(to_unsigned( 33,8)),
			1096 => std_logic_vector(to_unsigned( 119,8)),
			1097 => std_logic_vector(to_unsigned( 156,8)),
			1098 => std_logic_vector(to_unsigned( 162,8)),
			1099 => std_logic_vector(to_unsigned( 87,8)),
			1100 => std_logic_vector(to_unsigned( 149,8)),
			1101 => std_logic_vector(to_unsigned( 117,8)),
			1102 => std_logic_vector(to_unsigned( 28,8)),
			1103 => std_logic_vector(to_unsigned( 20,8)),
			1104 => std_logic_vector(to_unsigned( 42,8)),
			1105 => std_logic_vector(to_unsigned( 177,8)),
			1106 => std_logic_vector(to_unsigned( 132,8)),
			1107 => std_logic_vector(to_unsigned( 4,8)),
			1108 => std_logic_vector(to_unsigned( 106,8)),
			1109 => std_logic_vector(to_unsigned( 110,8)),
			1110 => std_logic_vector(to_unsigned( 248,8)),
			1111 => std_logic_vector(to_unsigned( 60,8)),
			1112 => std_logic_vector(to_unsigned( 154,8)),
			1113 => std_logic_vector(to_unsigned( 124,8)),
			1114 => std_logic_vector(to_unsigned( 30,8)),
			1115 => std_logic_vector(to_unsigned( 42,8)),
			1116 => std_logic_vector(to_unsigned( 165,8)),
			1117 => std_logic_vector(to_unsigned( 107,8)),
			1118 => std_logic_vector(to_unsigned( 217,8)),
			1119 => std_logic_vector(to_unsigned( 14,8)),
			1120 => std_logic_vector(to_unsigned( 19,8)),
			1121 => std_logic_vector(to_unsigned( 212,8)),
			1122 => std_logic_vector(to_unsigned( 185,8)),
			1123 => std_logic_vector(to_unsigned( 182,8)),
			1124 => std_logic_vector(to_unsigned( 56,8)),
			1125 => std_logic_vector(to_unsigned( 115,8)),
			1126 => std_logic_vector(to_unsigned( 123,8)),
			1127 => std_logic_vector(to_unsigned( 167,8)),
			1128 => std_logic_vector(to_unsigned( 241,8)),
			1129 => std_logic_vector(to_unsigned( 4,8)),
			1130 => std_logic_vector(to_unsigned( 18,8)),
			1131 => std_logic_vector(to_unsigned( 55,8)),
			1132 => std_logic_vector(to_unsigned( 24,8)),
			1133 => std_logic_vector(to_unsigned( 110,8)),
			1134 => std_logic_vector(to_unsigned( 42,8)),
			1135 => std_logic_vector(to_unsigned( 234,8)),
			1136 => std_logic_vector(to_unsigned( 136,8)),
			1137 => std_logic_vector(to_unsigned( 166,8)),
			1138 => std_logic_vector(to_unsigned( 67,8)),
			1139 => std_logic_vector(to_unsigned( 35,8)),
			1140 => std_logic_vector(to_unsigned( 1,8)),
			1141 => std_logic_vector(to_unsigned( 9,8)),
			1142 => std_logic_vector(to_unsigned( 15,8)),
			1143 => std_logic_vector(to_unsigned( 46,8)),
			1144 => std_logic_vector(to_unsigned( 196,8)),
			1145 => std_logic_vector(to_unsigned( 2,8)),
			1146 => std_logic_vector(to_unsigned( 93,8)),
			1147 => std_logic_vector(to_unsigned( 25,8)),
			1148 => std_logic_vector(to_unsigned( 140,8)),
			1149 => std_logic_vector(to_unsigned( 127,8)),
			1150 => std_logic_vector(to_unsigned( 121,8)),
			1151 => std_logic_vector(to_unsigned( 99,8)),
			1152 => std_logic_vector(to_unsigned( 206,8)),
			1153 => std_logic_vector(to_unsigned( 135,8)),
			1154 => std_logic_vector(to_unsigned( 160,8)),
			1155 => std_logic_vector(to_unsigned( 224,8)),
			1156 => std_logic_vector(to_unsigned( 255,8)),
			1157 => std_logic_vector(to_unsigned( 93,8)),
			1158 => std_logic_vector(to_unsigned( 215,8)),
			1159 => std_logic_vector(to_unsigned( 205,8)),
			1160 => std_logic_vector(to_unsigned( 228,8)),
			1161 => std_logic_vector(to_unsigned( 220,8)),
			1162 => std_logic_vector(to_unsigned( 87,8)),
			1163 => std_logic_vector(to_unsigned( 176,8)),
			1164 => std_logic_vector(to_unsigned( 93,8)),
			1165 => std_logic_vector(to_unsigned( 113,8)),
			1166 => std_logic_vector(to_unsigned( 208,8)),
			1167 => std_logic_vector(to_unsigned( 204,8)),
			1168 => std_logic_vector(to_unsigned( 190,8)),
			1169 => std_logic_vector(to_unsigned( 136,8)),
			1170 => std_logic_vector(to_unsigned( 108,8)),
			1171 => std_logic_vector(to_unsigned( 219,8)),
			1172 => std_logic_vector(to_unsigned( 93,8)),
			1173 => std_logic_vector(to_unsigned( 66,8)),
			1174 => std_logic_vector(to_unsigned( 115,8)),
			1175 => std_logic_vector(to_unsigned( 171,8)),
			1176 => std_logic_vector(to_unsigned( 165,8)),
			1177 => std_logic_vector(to_unsigned( 143,8)),
			1178 => std_logic_vector(to_unsigned( 31,8)),
			1179 => std_logic_vector(to_unsigned( 116,8)),
			1180 => std_logic_vector(to_unsigned( 167,8)),
			1181 => std_logic_vector(to_unsigned( 56,8)),
			1182 => std_logic_vector(to_unsigned( 231,8)),
			1183 => std_logic_vector(to_unsigned( 32,8)),
			1184 => std_logic_vector(to_unsigned( 238,8)),
			1185 => std_logic_vector(to_unsigned( 205,8)),
			1186 => std_logic_vector(to_unsigned( 55,8)),
			1187 => std_logic_vector(to_unsigned( 48,8)),
			1188 => std_logic_vector(to_unsigned( 147,8)),
			1189 => std_logic_vector(to_unsigned( 65,8)),
			1190 => std_logic_vector(to_unsigned( 224,8)),
			1191 => std_logic_vector(to_unsigned( 185,8)),
			1192 => std_logic_vector(to_unsigned( 243,8)),
			1193 => std_logic_vector(to_unsigned( 189,8)),
			1194 => std_logic_vector(to_unsigned( 163,8)),
			1195 => std_logic_vector(to_unsigned( 164,8)),
			1196 => std_logic_vector(to_unsigned( 154,8)),
			1197 => std_logic_vector(to_unsigned( 199,8)),
			1198 => std_logic_vector(to_unsigned( 98,8)),
			1199 => std_logic_vector(to_unsigned( 158,8)),
			1200 => std_logic_vector(to_unsigned( 176,8)),
			1201 => std_logic_vector(to_unsigned( 154,8)),
			1202 => std_logic_vector(to_unsigned( 183,8)),
			1203 => std_logic_vector(to_unsigned( 55,8)),
			1204 => std_logic_vector(to_unsigned( 210,8)),
			1205 => std_logic_vector(to_unsigned( 241,8)),
			1206 => std_logic_vector(to_unsigned( 14,8)),
			1207 => std_logic_vector(to_unsigned( 228,8)),
			1208 => std_logic_vector(to_unsigned( 46,8)),
			1209 => std_logic_vector(to_unsigned( 59,8)),
			1210 => std_logic_vector(to_unsigned( 17,8)),
			1211 => std_logic_vector(to_unsigned( 48,8)),
			1212 => std_logic_vector(to_unsigned( 211,8)),
			1213 => std_logic_vector(to_unsigned( 28,8)),
			1214 => std_logic_vector(to_unsigned( 33,8)),
			1215 => std_logic_vector(to_unsigned( 175,8)),
			1216 => std_logic_vector(to_unsigned( 145,8)),
			1217 => std_logic_vector(to_unsigned( 53,8)),
			1218 => std_logic_vector(to_unsigned( 231,8)),
			1219 => std_logic_vector(to_unsigned( 152,8)),
			1220 => std_logic_vector(to_unsigned( 39,8)),
			1221 => std_logic_vector(to_unsigned( 203,8)),
			1222 => std_logic_vector(to_unsigned( 73,8)),
			1223 => std_logic_vector(to_unsigned( 55,8)),
			1224 => std_logic_vector(to_unsigned( 165,8)),
			1225 => std_logic_vector(to_unsigned( 201,8)),
			1226 => std_logic_vector(to_unsigned( 209,8)),
			1227 => std_logic_vector(to_unsigned( 225,8)),
			1228 => std_logic_vector(to_unsigned( 130,8)),
			1229 => std_logic_vector(to_unsigned( 0,8)),
			1230 => std_logic_vector(to_unsigned( 107,8)),
			1231 => std_logic_vector(to_unsigned( 144,8)),
			1232 => std_logic_vector(to_unsigned( 133,8)),
			1233 => std_logic_vector(to_unsigned( 89,8)),
			1234 => std_logic_vector(to_unsigned( 137,8)),
			1235 => std_logic_vector(to_unsigned( 247,8)),
			1236 => std_logic_vector(to_unsigned( 158,8)),
			1237 => std_logic_vector(to_unsigned( 143,8)),
			1238 => std_logic_vector(to_unsigned( 108,8)),
			1239 => std_logic_vector(to_unsigned( 113,8)),
			1240 => std_logic_vector(to_unsigned( 239,8)),
			1241 => std_logic_vector(to_unsigned( 51,8)),
			1242 => std_logic_vector(to_unsigned( 186,8)),
			1243 => std_logic_vector(to_unsigned( 35,8)),
			1244 => std_logic_vector(to_unsigned( 39,8)),
			1245 => std_logic_vector(to_unsigned( 184,8)),
			1246 => std_logic_vector(to_unsigned( 133,8)),
			1247 => std_logic_vector(to_unsigned( 37,8)),
			1248 => std_logic_vector(to_unsigned( 250,8)),
			1249 => std_logic_vector(to_unsigned( 78,8)),
			1250 => std_logic_vector(to_unsigned( 230,8)),
			1251 => std_logic_vector(to_unsigned( 173,8)),
			1252 => std_logic_vector(to_unsigned( 141,8)),
			1253 => std_logic_vector(to_unsigned( 175,8)),
			1254 => std_logic_vector(to_unsigned( 4,8)),
			1255 => std_logic_vector(to_unsigned( 19,8)),
			1256 => std_logic_vector(to_unsigned( 104,8)),
			1257 => std_logic_vector(to_unsigned( 145,8)),
			1258 => std_logic_vector(to_unsigned( 184,8)),
			1259 => std_logic_vector(to_unsigned( 220,8)),
			1260 => std_logic_vector(to_unsigned( 146,8)),
			1261 => std_logic_vector(to_unsigned( 158,8)),
			1262 => std_logic_vector(to_unsigned( 141,8)),
			1263 => std_logic_vector(to_unsigned( 144,8)),
			1264 => std_logic_vector(to_unsigned( 191,8)),
			1265 => std_logic_vector(to_unsigned( 118,8)),
			1266 => std_logic_vector(to_unsigned( 36,8)),
			1267 => std_logic_vector(to_unsigned( 130,8)),
			1268 => std_logic_vector(to_unsigned( 76,8)),
			1269 => std_logic_vector(to_unsigned( 69,8)),
			1270 => std_logic_vector(to_unsigned( 184,8)),
			1271 => std_logic_vector(to_unsigned( 46,8)),
			1272 => std_logic_vector(to_unsigned( 146,8)),
			1273 => std_logic_vector(to_unsigned( 14,8)),
			1274 => std_logic_vector(to_unsigned( 192,8)),
			1275 => std_logic_vector(to_unsigned( 56,8)),
			1276 => std_logic_vector(to_unsigned( 128,8)),
			1277 => std_logic_vector(to_unsigned( 150,8)),
			1278 => std_logic_vector(to_unsigned( 201,8)),
			1279 => std_logic_vector(to_unsigned( 243,8)),
			1280 => std_logic_vector(to_unsigned( 85,8)),
			1281 => std_logic_vector(to_unsigned( 40,8)),
			1282 => std_logic_vector(to_unsigned( 199,8)),
			1283 => std_logic_vector(to_unsigned( 132,8)),
			1284 => std_logic_vector(to_unsigned( 175,8)),
			1285 => std_logic_vector(to_unsigned( 195,8)),
			1286 => std_logic_vector(to_unsigned( 255,8)),
			1287 => std_logic_vector(to_unsigned( 197,8)),
			1288 => std_logic_vector(to_unsigned( 236,8)),
			1289 => std_logic_vector(to_unsigned( 29,8)),
			1290 => std_logic_vector(to_unsigned( 70,8)),
			1291 => std_logic_vector(to_unsigned( 20,8)),
			1292 => std_logic_vector(to_unsigned( 75,8)),
			1293 => std_logic_vector(to_unsigned( 29,8)),
			1294 => std_logic_vector(to_unsigned( 163,8)),
			1295 => std_logic_vector(to_unsigned( 255,8)),
			1296 => std_logic_vector(to_unsigned( 155,8)),
			1297 => std_logic_vector(to_unsigned( 134,8)),
			1298 => std_logic_vector(to_unsigned( 89,8)),
			1299 => std_logic_vector(to_unsigned( 35,8)),
			1300 => std_logic_vector(to_unsigned( 98,8)),
			1301 => std_logic_vector(to_unsigned( 225,8)),
			1302 => std_logic_vector(to_unsigned( 190,8)),
			1303 => std_logic_vector(to_unsigned( 187,8)),
			1304 => std_logic_vector(to_unsigned( 111,8)),
			1305 => std_logic_vector(to_unsigned( 226,8)),
			1306 => std_logic_vector(to_unsigned( 93,8)),
			1307 => std_logic_vector(to_unsigned( 60,8)),
			1308 => std_logic_vector(to_unsigned( 175,8)),
			1309 => std_logic_vector(to_unsigned( 139,8)),
			1310 => std_logic_vector(to_unsigned( 181,8)),
			1311 => std_logic_vector(to_unsigned( 100,8)),
			1312 => std_logic_vector(to_unsigned( 207,8)),
			1313 => std_logic_vector(to_unsigned( 77,8)),
			1314 => std_logic_vector(to_unsigned( 11,8)),
			1315 => std_logic_vector(to_unsigned( 185,8)),
			1316 => std_logic_vector(to_unsigned( 234,8)),
			1317 => std_logic_vector(to_unsigned( 65,8)),
			1318 => std_logic_vector(to_unsigned( 179,8)),
			1319 => std_logic_vector(to_unsigned( 184,8)),
			1320 => std_logic_vector(to_unsigned( 245,8)),
			1321 => std_logic_vector(to_unsigned( 45,8)),
			1322 => std_logic_vector(to_unsigned( 244,8)),
			1323 => std_logic_vector(to_unsigned( 1,8)),
			1324 => std_logic_vector(to_unsigned( 238,8)),
			1325 => std_logic_vector(to_unsigned( 8,8)),
			1326 => std_logic_vector(to_unsigned( 219,8)),
			1327 => std_logic_vector(to_unsigned( 213,8)),
			1328 => std_logic_vector(to_unsigned( 3,8)),
			1329 => std_logic_vector(to_unsigned( 32,8)),
			1330 => std_logic_vector(to_unsigned( 55,8)),
			1331 => std_logic_vector(to_unsigned( 226,8)),
			1332 => std_logic_vector(to_unsigned( 37,8)),
			1333 => std_logic_vector(to_unsigned( 24,8)),
			1334 => std_logic_vector(to_unsigned( 139,8)),
			1335 => std_logic_vector(to_unsigned( 138,8)),
			1336 => std_logic_vector(to_unsigned( 59,8)),
			1337 => std_logic_vector(to_unsigned( 226,8)),
			1338 => std_logic_vector(to_unsigned( 224,8)),
			1339 => std_logic_vector(to_unsigned( 123,8)),
			1340 => std_logic_vector(to_unsigned( 27,8)),
			1341 => std_logic_vector(to_unsigned( 135,8)),
			1342 => std_logic_vector(to_unsigned( 87,8)),
			1343 => std_logic_vector(to_unsigned( 27,8)),
			1344 => std_logic_vector(to_unsigned( 11,8)),
			1345 => std_logic_vector(to_unsigned( 99,8)),
			1346 => std_logic_vector(to_unsigned( 225,8)),
			1347 => std_logic_vector(to_unsigned( 132,8)),
			1348 => std_logic_vector(to_unsigned( 192,8)),
			1349 => std_logic_vector(to_unsigned( 177,8)),
			1350 => std_logic_vector(to_unsigned( 33,8)),
			1351 => std_logic_vector(to_unsigned( 209,8)),
			1352 => std_logic_vector(to_unsigned( 220,8)),
			1353 => std_logic_vector(to_unsigned( 216,8)),
			1354 => std_logic_vector(to_unsigned( 79,8)),
			1355 => std_logic_vector(to_unsigned( 26,8)),
			1356 => std_logic_vector(to_unsigned( 132,8)),
			1357 => std_logic_vector(to_unsigned( 47,8)),
			1358 => std_logic_vector(to_unsigned( 134,8)),
			1359 => std_logic_vector(to_unsigned( 252,8)),
			1360 => std_logic_vector(to_unsigned( 200,8)),
			1361 => std_logic_vector(to_unsigned( 56,8)),
			1362 => std_logic_vector(to_unsigned( 233,8)),
			1363 => std_logic_vector(to_unsigned( 66,8)),
			1364 => std_logic_vector(to_unsigned( 189,8)),
			1365 => std_logic_vector(to_unsigned( 224,8)),
			1366 => std_logic_vector(to_unsigned( 127,8)),
			1367 => std_logic_vector(to_unsigned( 32,8)),
			1368 => std_logic_vector(to_unsigned( 128,8)),
			1369 => std_logic_vector(to_unsigned( 132,8)),
			1370 => std_logic_vector(to_unsigned( 103,8)),
			1371 => std_logic_vector(to_unsigned( 57,8)),
			1372 => std_logic_vector(to_unsigned( 103,8)),
			1373 => std_logic_vector(to_unsigned( 197,8)),
			1374 => std_logic_vector(to_unsigned( 15,8)),
			1375 => std_logic_vector(to_unsigned( 60,8)),
			1376 => std_logic_vector(to_unsigned( 250,8)),
			1377 => std_logic_vector(to_unsigned( 246,8)),
			1378 => std_logic_vector(to_unsigned( 198,8)),
			1379 => std_logic_vector(to_unsigned( 158,8)),
			1380 => std_logic_vector(to_unsigned( 24,8)),
			1381 => std_logic_vector(to_unsigned( 124,8)),
			1382 => std_logic_vector(to_unsigned( 218,8)),
			1383 => std_logic_vector(to_unsigned( 32,8)),
			1384 => std_logic_vector(to_unsigned( 153,8)),
			1385 => std_logic_vector(to_unsigned( 241,8)),
			1386 => std_logic_vector(to_unsigned( 37,8)),
			1387 => std_logic_vector(to_unsigned( 5,8)),
			1388 => std_logic_vector(to_unsigned( 252,8)),
			1389 => std_logic_vector(to_unsigned( 136,8)),
			1390 => std_logic_vector(to_unsigned( 246,8)),
			1391 => std_logic_vector(to_unsigned( 192,8)),
			1392 => std_logic_vector(to_unsigned( 194,8)),
			1393 => std_logic_vector(to_unsigned( 83,8)),
			1394 => std_logic_vector(to_unsigned( 4,8)),
			1395 => std_logic_vector(to_unsigned( 148,8)),
			1396 => std_logic_vector(to_unsigned( 223,8)),
			1397 => std_logic_vector(to_unsigned( 49,8)),
			1398 => std_logic_vector(to_unsigned( 143,8)),
			1399 => std_logic_vector(to_unsigned( 78,8)),
			1400 => std_logic_vector(to_unsigned( 107,8)),
			1401 => std_logic_vector(to_unsigned( 215,8)),
			1402 => std_logic_vector(to_unsigned( 118,8)),
			1403 => std_logic_vector(to_unsigned( 211,8)),
			1404 => std_logic_vector(to_unsigned( 177,8)),
			1405 => std_logic_vector(to_unsigned( 90,8)),
			1406 => std_logic_vector(to_unsigned( 162,8)),
			1407 => std_logic_vector(to_unsigned( 118,8)),
			1408 => std_logic_vector(to_unsigned( 116,8)),
			1409 => std_logic_vector(to_unsigned( 174,8)),
			1410 => std_logic_vector(to_unsigned( 47,8)),
			1411 => std_logic_vector(to_unsigned( 40,8)),
			1412 => std_logic_vector(to_unsigned( 40,8)),
			1413 => std_logic_vector(to_unsigned( 202,8)),
			1414 => std_logic_vector(to_unsigned( 14,8)),
			1415 => std_logic_vector(to_unsigned( 77,8)),
			1416 => std_logic_vector(to_unsigned( 70,8)),
			1417 => std_logic_vector(to_unsigned( 62,8)),
			1418 => std_logic_vector(to_unsigned( 101,8)),
			1419 => std_logic_vector(to_unsigned( 193,8)),
			1420 => std_logic_vector(to_unsigned( 158,8)),
			1421 => std_logic_vector(to_unsigned( 57,8)),
			1422 => std_logic_vector(to_unsigned( 144,8)),
			1423 => std_logic_vector(to_unsigned( 121,8)),
			1424 => std_logic_vector(to_unsigned( 118,8)),
			1425 => std_logic_vector(to_unsigned( 122,8)),
			1426 => std_logic_vector(to_unsigned( 245,8)),
			1427 => std_logic_vector(to_unsigned( 189,8)),
			1428 => std_logic_vector(to_unsigned( 243,8)),
			1429 => std_logic_vector(to_unsigned( 124,8)),
			1430 => std_logic_vector(to_unsigned( 27,8)),
			1431 => std_logic_vector(to_unsigned( 127,8)),
			1432 => std_logic_vector(to_unsigned( 73,8)),
			1433 => std_logic_vector(to_unsigned( 225,8)),
			1434 => std_logic_vector(to_unsigned( 154,8)),
			1435 => std_logic_vector(to_unsigned( 227,8)),
			1436 => std_logic_vector(to_unsigned( 99,8)),
			1437 => std_logic_vector(to_unsigned( 100,8)),
			1438 => std_logic_vector(to_unsigned( 237,8)),
			1439 => std_logic_vector(to_unsigned( 168,8)),
			1440 => std_logic_vector(to_unsigned( 2,8)),
			1441 => std_logic_vector(to_unsigned( 171,8)),
			1442 => std_logic_vector(to_unsigned( 235,8)),
			1443 => std_logic_vector(to_unsigned( 63,8)),
			1444 => std_logic_vector(to_unsigned( 91,8)),
			1445 => std_logic_vector(to_unsigned( 30,8)),
			1446 => std_logic_vector(to_unsigned( 74,8)),
			1447 => std_logic_vector(to_unsigned( 17,8)),
			1448 => std_logic_vector(to_unsigned( 84,8)),
			1449 => std_logic_vector(to_unsigned( 214,8)),
			1450 => std_logic_vector(to_unsigned( 151,8)),
			1451 => std_logic_vector(to_unsigned( 197,8)),
			1452 => std_logic_vector(to_unsigned( 94,8)),
			1453 => std_logic_vector(to_unsigned( 56,8)),
			1454 => std_logic_vector(to_unsigned( 9,8)),
			1455 => std_logic_vector(to_unsigned( 237,8)),
			1456 => std_logic_vector(to_unsigned( 111,8)),
			1457 => std_logic_vector(to_unsigned( 176,8)),
			1458 => std_logic_vector(to_unsigned( 196,8)),
			1459 => std_logic_vector(to_unsigned( 234,8)),
			1460 => std_logic_vector(to_unsigned( 228,8)),
			1461 => std_logic_vector(to_unsigned( 34,8)),
			1462 => std_logic_vector(to_unsigned( 89,8)),
			1463 => std_logic_vector(to_unsigned( 188,8)),
			1464 => std_logic_vector(to_unsigned( 168,8)),
			1465 => std_logic_vector(to_unsigned( 180,8)),
			1466 => std_logic_vector(to_unsigned( 49,8)),
			1467 => std_logic_vector(to_unsigned( 166,8)),
			1468 => std_logic_vector(to_unsigned( 246,8)),
			1469 => std_logic_vector(to_unsigned( 77,8)),
			1470 => std_logic_vector(to_unsigned( 28,8)),
			1471 => std_logic_vector(to_unsigned( 81,8)),
			1472 => std_logic_vector(to_unsigned( 166,8)),
			1473 => std_logic_vector(to_unsigned( 87,8)),
			1474 => std_logic_vector(to_unsigned( 113,8)),
			1475 => std_logic_vector(to_unsigned( 254,8)),
			1476 => std_logic_vector(to_unsigned( 219,8)),
			1477 => std_logic_vector(to_unsigned( 138,8)),
			1478 => std_logic_vector(to_unsigned( 101,8)),
			1479 => std_logic_vector(to_unsigned( 23,8)),
			1480 => std_logic_vector(to_unsigned( 249,8)),
			1481 => std_logic_vector(to_unsigned( 50,8)),
			1482 => std_logic_vector(to_unsigned( 28,8)),
			1483 => std_logic_vector(to_unsigned( 54,8)),
			1484 => std_logic_vector(to_unsigned( 237,8)),
			1485 => std_logic_vector(to_unsigned( 235,8)),
			1486 => std_logic_vector(to_unsigned( 152,8)),
			1487 => std_logic_vector(to_unsigned( 60,8)),
			1488 => std_logic_vector(to_unsigned( 69,8)),
			1489 => std_logic_vector(to_unsigned( 205,8)),
			1490 => std_logic_vector(to_unsigned( 70,8)),
			1491 => std_logic_vector(to_unsigned( 208,8)),
			1492 => std_logic_vector(to_unsigned( 57,8)),
			1493 => std_logic_vector(to_unsigned( 21,8)),
			1494 => std_logic_vector(to_unsigned( 223,8)),
			1495 => std_logic_vector(to_unsigned( 99,8)),
			1496 => std_logic_vector(to_unsigned( 137,8)),
			1497 => std_logic_vector(to_unsigned( 234,8)),
			1498 => std_logic_vector(to_unsigned( 55,8)),
			1499 => std_logic_vector(to_unsigned( 5,8)),
			1500 => std_logic_vector(to_unsigned( 167,8)),
			1501 => std_logic_vector(to_unsigned( 250,8)),
			1502 => std_logic_vector(to_unsigned( 29,8)),
			1503 => std_logic_vector(to_unsigned( 87,8)),
			1504 => std_logic_vector(to_unsigned( 158,8)),
			1505 => std_logic_vector(to_unsigned( 152,8)),
			1506 => std_logic_vector(to_unsigned( 64,8)),
			1507 => std_logic_vector(to_unsigned( 216,8)),
			1508 => std_logic_vector(to_unsigned( 82,8)),
			1509 => std_logic_vector(to_unsigned( 120,8)),
			1510 => std_logic_vector(to_unsigned( 23,8)),
			1511 => std_logic_vector(to_unsigned( 44,8)),
			1512 => std_logic_vector(to_unsigned( 212,8)),
			1513 => std_logic_vector(to_unsigned( 253,8)),
			1514 => std_logic_vector(to_unsigned( 16,8)),
			1515 => std_logic_vector(to_unsigned( 195,8)),
			1516 => std_logic_vector(to_unsigned( 236,8)),
			1517 => std_logic_vector(to_unsigned( 148,8)),
			1518 => std_logic_vector(to_unsigned( 48,8)),
			1519 => std_logic_vector(to_unsigned( 252,8)),
			1520 => std_logic_vector(to_unsigned( 56,8)),
			1521 => std_logic_vector(to_unsigned( 69,8)),
			1522 => std_logic_vector(to_unsigned( 158,8)),
			1523 => std_logic_vector(to_unsigned( 248,8)),
			1524 => std_logic_vector(to_unsigned( 102,8)),
			1525 => std_logic_vector(to_unsigned( 55,8)),
			1526 => std_logic_vector(to_unsigned( 16,8)),
			1527 => std_logic_vector(to_unsigned( 140,8)),
			1528 => std_logic_vector(to_unsigned( 140,8)),
			1529 => std_logic_vector(to_unsigned( 185,8)),
			1530 => std_logic_vector(to_unsigned( 169,8)),
			1531 => std_logic_vector(to_unsigned( 235,8)),
			1532 => std_logic_vector(to_unsigned( 134,8)),
			1533 => std_logic_vector(to_unsigned( 143,8)),
			1534 => std_logic_vector(to_unsigned( 165,8)),
			1535 => std_logic_vector(to_unsigned( 34,8)),
			1536 => std_logic_vector(to_unsigned( 92,8)),
			1537 => std_logic_vector(to_unsigned( 170,8)),
			1538 => std_logic_vector(to_unsigned( 180,8)),
			1539 => std_logic_vector(to_unsigned( 89,8)),
			1540 => std_logic_vector(to_unsigned( 172,8)),
			1541 => std_logic_vector(to_unsigned( 82,8)),
			1542 => std_logic_vector(to_unsigned( 222,8)),
			1543 => std_logic_vector(to_unsigned( 169,8)),
			1544 => std_logic_vector(to_unsigned( 118,8)),
			1545 => std_logic_vector(to_unsigned( 193,8)),
			1546 => std_logic_vector(to_unsigned( 148,8)),
			1547 => std_logic_vector(to_unsigned( 229,8)),
			1548 => std_logic_vector(to_unsigned( 188,8)),
			1549 => std_logic_vector(to_unsigned( 207,8)),
			1550 => std_logic_vector(to_unsigned( 228,8)),
			1551 => std_logic_vector(to_unsigned( 8,8)),
			1552 => std_logic_vector(to_unsigned( 111,8)),
			1553 => std_logic_vector(to_unsigned( 107,8)),
			1554 => std_logic_vector(to_unsigned( 88,8)),
			1555 => std_logic_vector(to_unsigned( 3,8)),
			1556 => std_logic_vector(to_unsigned( 211,8)),
			1557 => std_logic_vector(to_unsigned( 122,8)),
			1558 => std_logic_vector(to_unsigned( 55,8)),
			1559 => std_logic_vector(to_unsigned( 182,8)),
			1560 => std_logic_vector(to_unsigned( 195,8)),
			1561 => std_logic_vector(to_unsigned( 136,8)),
			1562 => std_logic_vector(to_unsigned( 229,8)),
			1563 => std_logic_vector(to_unsigned( 206,8)),
			1564 => std_logic_vector(to_unsigned( 79,8)),
			1565 => std_logic_vector(to_unsigned( 102,8)),
			1566 => std_logic_vector(to_unsigned( 241,8)),
			1567 => std_logic_vector(to_unsigned( 197,8)),
			1568 => std_logic_vector(to_unsigned( 214,8)),
			1569 => std_logic_vector(to_unsigned( 137,8)),
			1570 => std_logic_vector(to_unsigned( 21,8)),
			1571 => std_logic_vector(to_unsigned( 42,8)),
			1572 => std_logic_vector(to_unsigned( 203,8)),
			1573 => std_logic_vector(to_unsigned( 58,8)),
			1574 => std_logic_vector(to_unsigned( 222,8)),
			1575 => std_logic_vector(to_unsigned( 17,8)),
			1576 => std_logic_vector(to_unsigned( 138,8)),
			1577 => std_logic_vector(to_unsigned( 123,8)),
			1578 => std_logic_vector(to_unsigned( 175,8)),
			1579 => std_logic_vector(to_unsigned( 36,8)),
			1580 => std_logic_vector(to_unsigned( 89,8)),
			1581 => std_logic_vector(to_unsigned( 253,8)),
			1582 => std_logic_vector(to_unsigned( 254,8)),
			1583 => std_logic_vector(to_unsigned( 250,8)),
			1584 => std_logic_vector(to_unsigned( 148,8)),
			1585 => std_logic_vector(to_unsigned( 60,8)),
			1586 => std_logic_vector(to_unsigned( 251,8)),
			1587 => std_logic_vector(to_unsigned( 105,8)),
			1588 => std_logic_vector(to_unsigned( 45,8)),
			1589 => std_logic_vector(to_unsigned( 160,8)),
			1590 => std_logic_vector(to_unsigned( 151,8)),
			1591 => std_logic_vector(to_unsigned( 161,8)),
			1592 => std_logic_vector(to_unsigned( 15,8)),
			1593 => std_logic_vector(to_unsigned( 180,8)),
			1594 => std_logic_vector(to_unsigned( 71,8)),
			1595 => std_logic_vector(to_unsigned( 5,8)),
			1596 => std_logic_vector(to_unsigned( 196,8)),
			1597 => std_logic_vector(to_unsigned( 133,8)),
			1598 => std_logic_vector(to_unsigned( 164,8)),
			1599 => std_logic_vector(to_unsigned( 201,8)),
			1600 => std_logic_vector(to_unsigned( 224,8)),
			1601 => std_logic_vector(to_unsigned( 51,8)),
			1602 => std_logic_vector(to_unsigned( 193,8)),
			1603 => std_logic_vector(to_unsigned( 122,8)),
			1604 => std_logic_vector(to_unsigned( 135,8)),
			1605 => std_logic_vector(to_unsigned( 104,8)),
			1606 => std_logic_vector(to_unsigned( 70,8)),
			1607 => std_logic_vector(to_unsigned( 48,8)),
			1608 => std_logic_vector(to_unsigned( 46,8)),
			1609 => std_logic_vector(to_unsigned( 26,8)),
			1610 => std_logic_vector(to_unsigned( 206,8)),
			1611 => std_logic_vector(to_unsigned( 183,8)),
			1612 => std_logic_vector(to_unsigned( 215,8)),
			1613 => std_logic_vector(to_unsigned( 187,8)),
			1614 => std_logic_vector(to_unsigned( 18,8)),
			1615 => std_logic_vector(to_unsigned( 113,8)),
			1616 => std_logic_vector(to_unsigned( 71,8)),
			1617 => std_logic_vector(to_unsigned( 160,8)),
			1618 => std_logic_vector(to_unsigned( 14,8)),
			1619 => std_logic_vector(to_unsigned( 137,8)),
			1620 => std_logic_vector(to_unsigned( 202,8)),
			1621 => std_logic_vector(to_unsigned( 95,8)),
			1622 => std_logic_vector(to_unsigned( 229,8)),
			1623 => std_logic_vector(to_unsigned( 91,8)),
			1624 => std_logic_vector(to_unsigned( 201,8)),
			1625 => std_logic_vector(to_unsigned( 42,8)),
			1626 => std_logic_vector(to_unsigned( 215,8)),
			1627 => std_logic_vector(to_unsigned( 151,8)),
			1628 => std_logic_vector(to_unsigned( 96,8)),
			1629 => std_logic_vector(to_unsigned( 55,8)),
			1630 => std_logic_vector(to_unsigned( 113,8)),
			1631 => std_logic_vector(to_unsigned( 29,8)),
			1632 => std_logic_vector(to_unsigned( 104,8)),
			1633 => std_logic_vector(to_unsigned( 140,8)),
			1634 => std_logic_vector(to_unsigned( 174,8)),
			1635 => std_logic_vector(to_unsigned( 165,8)),
			1636 => std_logic_vector(to_unsigned( 37,8)),
			1637 => std_logic_vector(to_unsigned( 178,8)),
			1638 => std_logic_vector(to_unsigned( 143,8)),
			1639 => std_logic_vector(to_unsigned( 185,8)),
			1640 => std_logic_vector(to_unsigned( 252,8)),
			1641 => std_logic_vector(to_unsigned( 174,8)),
			1642 => std_logic_vector(to_unsigned( 253,8)),
			1643 => std_logic_vector(to_unsigned( 134,8)),
			1644 => std_logic_vector(to_unsigned( 77,8)),
			1645 => std_logic_vector(to_unsigned( 99,8)),
			1646 => std_logic_vector(to_unsigned( 39,8)),
			1647 => std_logic_vector(to_unsigned( 136,8)),
			1648 => std_logic_vector(to_unsigned( 143,8)),
			1649 => std_logic_vector(to_unsigned( 128,8)),
			1650 => std_logic_vector(to_unsigned( 90,8)),
			1651 => std_logic_vector(to_unsigned( 188,8)),
			1652 => std_logic_vector(to_unsigned( 69,8)),
			1653 => std_logic_vector(to_unsigned( 88,8)),
			1654 => std_logic_vector(to_unsigned( 108,8)),
			1655 => std_logic_vector(to_unsigned( 53,8)),
			1656 => std_logic_vector(to_unsigned( 22,8)),
			1657 => std_logic_vector(to_unsigned( 216,8)),
			1658 => std_logic_vector(to_unsigned( 63,8)),
			1659 => std_logic_vector(to_unsigned( 207,8)),
			1660 => std_logic_vector(to_unsigned( 27,8)),
			1661 => std_logic_vector(to_unsigned( 238,8)),
			1662 => std_logic_vector(to_unsigned( 179,8)),
			1663 => std_logic_vector(to_unsigned( 56,8)),
			1664 => std_logic_vector(to_unsigned( 85,8)),
			1665 => std_logic_vector(to_unsigned( 71,8)),
			1666 => std_logic_vector(to_unsigned( 73,8)),
			1667 => std_logic_vector(to_unsigned( 102,8)),
			1668 => std_logic_vector(to_unsigned( 162,8)),
			1669 => std_logic_vector(to_unsigned( 3,8)),
			1670 => std_logic_vector(to_unsigned( 90,8)),
			1671 => std_logic_vector(to_unsigned( 81,8)),
			1672 => std_logic_vector(to_unsigned( 74,8)),
			1673 => std_logic_vector(to_unsigned( 122,8)),
			1674 => std_logic_vector(to_unsigned( 54,8)),
			1675 => std_logic_vector(to_unsigned( 209,8)),
			1676 => std_logic_vector(to_unsigned( 18,8)),
			1677 => std_logic_vector(to_unsigned( 223,8)),
			1678 => std_logic_vector(to_unsigned( 41,8)),
			1679 => std_logic_vector(to_unsigned( 75,8)),
			1680 => std_logic_vector(to_unsigned( 36,8)),
			1681 => std_logic_vector(to_unsigned( 38,8)),
			1682 => std_logic_vector(to_unsigned( 196,8)),
			1683 => std_logic_vector(to_unsigned( 62,8)),
			1684 => std_logic_vector(to_unsigned( 108,8)),
			1685 => std_logic_vector(to_unsigned( 108,8)),
			1686 => std_logic_vector(to_unsigned( 224,8)),
			1687 => std_logic_vector(to_unsigned( 0,8)),
			1688 => std_logic_vector(to_unsigned( 227,8)),
			1689 => std_logic_vector(to_unsigned( 187,8)),
			1690 => std_logic_vector(to_unsigned( 224,8)),
			1691 => std_logic_vector(to_unsigned( 147,8)),
			1692 => std_logic_vector(to_unsigned( 177,8)),
			1693 => std_logic_vector(to_unsigned( 140,8)),
			1694 => std_logic_vector(to_unsigned( 36,8)),
			1695 => std_logic_vector(to_unsigned( 113,8)),
			1696 => std_logic_vector(to_unsigned( 140,8)),
			1697 => std_logic_vector(to_unsigned( 241,8)),
			1698 => std_logic_vector(to_unsigned( 21,8)),
			1699 => std_logic_vector(to_unsigned( 135,8)),
			1700 => std_logic_vector(to_unsigned( 17,8)),
			1701 => std_logic_vector(to_unsigned( 98,8)),
			1702 => std_logic_vector(to_unsigned( 103,8)),
			1703 => std_logic_vector(to_unsigned( 21,8)),
			1704 => std_logic_vector(to_unsigned( 46,8)),
			1705 => std_logic_vector(to_unsigned( 177,8)),
			1706 => std_logic_vector(to_unsigned( 89,8)),
			1707 => std_logic_vector(to_unsigned( 152,8)),
			1708 => std_logic_vector(to_unsigned( 81,8)),
			1709 => std_logic_vector(to_unsigned( 136,8)),
			1710 => std_logic_vector(to_unsigned( 124,8)),
			1711 => std_logic_vector(to_unsigned( 211,8)),
			1712 => std_logic_vector(to_unsigned( 139,8)),
			1713 => std_logic_vector(to_unsigned( 147,8)),
			1714 => std_logic_vector(to_unsigned( 14,8)),
			1715 => std_logic_vector(to_unsigned( 75,8)),
			1716 => std_logic_vector(to_unsigned( 221,8)),
			1717 => std_logic_vector(to_unsigned( 179,8)),
			1718 => std_logic_vector(to_unsigned( 204,8)),
			1719 => std_logic_vector(to_unsigned( 95,8)),
			1720 => std_logic_vector(to_unsigned( 121,8)),
			1721 => std_logic_vector(to_unsigned( 7,8)),
			1722 => std_logic_vector(to_unsigned( 190,8)),
			1723 => std_logic_vector(to_unsigned( 130,8)),
			1724 => std_logic_vector(to_unsigned( 198,8)),
			1725 => std_logic_vector(to_unsigned( 142,8)),
			1726 => std_logic_vector(to_unsigned( 141,8)),
			1727 => std_logic_vector(to_unsigned( 184,8)),
			1728 => std_logic_vector(to_unsigned( 159,8)),
			1729 => std_logic_vector(to_unsigned( 215,8)),
			1730 => std_logic_vector(to_unsigned( 7,8)),
			1731 => std_logic_vector(to_unsigned( 225,8)),
			1732 => std_logic_vector(to_unsigned( 104,8)),
			1733 => std_logic_vector(to_unsigned( 91,8)),
			1734 => std_logic_vector(to_unsigned( 232,8)),
			1735 => std_logic_vector(to_unsigned( 32,8)),
			1736 => std_logic_vector(to_unsigned( 207,8)),
			1737 => std_logic_vector(to_unsigned( 125,8)),
			1738 => std_logic_vector(to_unsigned( 242,8)),
			1739 => std_logic_vector(to_unsigned( 242,8)),
			1740 => std_logic_vector(to_unsigned( 0,8)),
			1741 => std_logic_vector(to_unsigned( 122,8)),
			1742 => std_logic_vector(to_unsigned( 192,8)),
			1743 => std_logic_vector(to_unsigned( 215,8)),
			1744 => std_logic_vector(to_unsigned( 108,8)),
			1745 => std_logic_vector(to_unsigned( 220,8)),
			1746 => std_logic_vector(to_unsigned( 254,8)),
			1747 => std_logic_vector(to_unsigned( 192,8)),
			1748 => std_logic_vector(to_unsigned( 162,8)),
			1749 => std_logic_vector(to_unsigned( 60,8)),
			1750 => std_logic_vector(to_unsigned( 188,8)),
			1751 => std_logic_vector(to_unsigned( 64,8)),
			1752 => std_logic_vector(to_unsigned( 72,8)),
			1753 => std_logic_vector(to_unsigned( 120,8)),
			1754 => std_logic_vector(to_unsigned( 230,8)),
			1755 => std_logic_vector(to_unsigned( 175,8)),
			1756 => std_logic_vector(to_unsigned( 196,8)),
			1757 => std_logic_vector(to_unsigned( 98,8)),
			1758 => std_logic_vector(to_unsigned( 232,8)),
			1759 => std_logic_vector(to_unsigned( 127,8)),
			1760 => std_logic_vector(to_unsigned( 81,8)),
			1761 => std_logic_vector(to_unsigned( 66,8)),
			1762 => std_logic_vector(to_unsigned( 105,8)),
			1763 => std_logic_vector(to_unsigned( 167,8)),
			1764 => std_logic_vector(to_unsigned( 192,8)),
			1765 => std_logic_vector(to_unsigned( 29,8)),
			1766 => std_logic_vector(to_unsigned( 246,8)),
			1767 => std_logic_vector(to_unsigned( 114,8)),
			1768 => std_logic_vector(to_unsigned( 25,8)),
			1769 => std_logic_vector(to_unsigned( 87,8)),
			1770 => std_logic_vector(to_unsigned( 123,8)),
			1771 => std_logic_vector(to_unsigned( 220,8)),
			1772 => std_logic_vector(to_unsigned( 102,8)),
			1773 => std_logic_vector(to_unsigned( 104,8)),
			1774 => std_logic_vector(to_unsigned( 54,8)),
			1775 => std_logic_vector(to_unsigned( 24,8)),
			1776 => std_logic_vector(to_unsigned( 87,8)),
			1777 => std_logic_vector(to_unsigned( 229,8)),
			1778 => std_logic_vector(to_unsigned( 178,8)),
			1779 => std_logic_vector(to_unsigned( 60,8)),
			1780 => std_logic_vector(to_unsigned( 226,8)),
			1781 => std_logic_vector(to_unsigned( 103,8)),
			1782 => std_logic_vector(to_unsigned( 71,8)),
			1783 => std_logic_vector(to_unsigned( 54,8)),
			1784 => std_logic_vector(to_unsigned( 76,8)),
			1785 => std_logic_vector(to_unsigned( 51,8)),
			1786 => std_logic_vector(to_unsigned( 118,8)),
			1787 => std_logic_vector(to_unsigned( 134,8)),
			1788 => std_logic_vector(to_unsigned( 20,8)),
			1789 => std_logic_vector(to_unsigned( 66,8)),
			1790 => std_logic_vector(to_unsigned( 85,8)),
			1791 => std_logic_vector(to_unsigned( 143,8)),
			1792 => std_logic_vector(to_unsigned( 251,8)),
			1793 => std_logic_vector(to_unsigned( 85,8)),
			1794 => std_logic_vector(to_unsigned( 197,8)),
			1795 => std_logic_vector(to_unsigned( 112,8)),
			1796 => std_logic_vector(to_unsigned( 100,8)),
			1797 => std_logic_vector(to_unsigned( 137,8)),
			1798 => std_logic_vector(to_unsigned( 50,8)),
			1799 => std_logic_vector(to_unsigned( 227,8)),
			1800 => std_logic_vector(to_unsigned( 176,8)),
			1801 => std_logic_vector(to_unsigned( 186,8)),
			1802 => std_logic_vector(to_unsigned( 78,8)),
			1803 => std_logic_vector(to_unsigned( 63,8)),
			1804 => std_logic_vector(to_unsigned( 238,8)),
			1805 => std_logic_vector(to_unsigned( 104,8)),
			1806 => std_logic_vector(to_unsigned( 140,8)),
			1807 => std_logic_vector(to_unsigned( 16,8)),
			1808 => std_logic_vector(to_unsigned( 208,8)),
			1809 => std_logic_vector(to_unsigned( 43,8)),
			1810 => std_logic_vector(to_unsigned( 117,8)),
			1811 => std_logic_vector(to_unsigned( 148,8)),
			1812 => std_logic_vector(to_unsigned( 28,8)),
			1813 => std_logic_vector(to_unsigned( 53,8)),
			1814 => std_logic_vector(to_unsigned( 83,8)),
			1815 => std_logic_vector(to_unsigned( 192,8)),
			1816 => std_logic_vector(to_unsigned( 226,8)),
			1817 => std_logic_vector(to_unsigned( 177,8)),
			1818 => std_logic_vector(to_unsigned( 77,8)),
			1819 => std_logic_vector(to_unsigned( 19,8)),
			1820 => std_logic_vector(to_unsigned( 200,8)),
			1821 => std_logic_vector(to_unsigned( 185,8)),
			1822 => std_logic_vector(to_unsigned( 149,8)),
			1823 => std_logic_vector(to_unsigned( 142,8)),
			1824 => std_logic_vector(to_unsigned( 57,8)),
			1825 => std_logic_vector(to_unsigned( 177,8)),
			1826 => std_logic_vector(to_unsigned( 19,8)),
			1827 => std_logic_vector(to_unsigned( 158,8)),
			1828 => std_logic_vector(to_unsigned( 245,8)),
			1829 => std_logic_vector(to_unsigned( 77,8)),
			1830 => std_logic_vector(to_unsigned( 161,8)),
			1831 => std_logic_vector(to_unsigned( 27,8)),
			1832 => std_logic_vector(to_unsigned( 222,8)),
			1833 => std_logic_vector(to_unsigned( 108,8)),
			1834 => std_logic_vector(to_unsigned( 74,8)),
			1835 => std_logic_vector(to_unsigned( 45,8)),
			1836 => std_logic_vector(to_unsigned( 66,8)),
			1837 => std_logic_vector(to_unsigned( 162,8)),
			1838 => std_logic_vector(to_unsigned( 111,8)),
			1839 => std_logic_vector(to_unsigned( 35,8)),
			1840 => std_logic_vector(to_unsigned( 118,8)),
			1841 => std_logic_vector(to_unsigned( 116,8)),
			1842 => std_logic_vector(to_unsigned( 139,8)),
			1843 => std_logic_vector(to_unsigned( 252,8)),
			1844 => std_logic_vector(to_unsigned( 66,8)),
			1845 => std_logic_vector(to_unsigned( 56,8)),
			1846 => std_logic_vector(to_unsigned( 2,8)),
			1847 => std_logic_vector(to_unsigned( 235,8)),
			1848 => std_logic_vector(to_unsigned( 70,8)),
			1849 => std_logic_vector(to_unsigned( 153,8)),
			1850 => std_logic_vector(to_unsigned( 35,8)),
			1851 => std_logic_vector(to_unsigned( 127,8)),
			1852 => std_logic_vector(to_unsigned( 224,8)),
			1853 => std_logic_vector(to_unsigned( 188,8)),
			1854 => std_logic_vector(to_unsigned( 251,8)),
			1855 => std_logic_vector(to_unsigned( 85,8)),
			1856 => std_logic_vector(to_unsigned( 125,8)),
			1857 => std_logic_vector(to_unsigned( 251,8)),
			1858 => std_logic_vector(to_unsigned( 27,8)),
			1859 => std_logic_vector(to_unsigned( 169,8)),
			1860 => std_logic_vector(to_unsigned( 97,8)),
			1861 => std_logic_vector(to_unsigned( 115,8)),
			1862 => std_logic_vector(to_unsigned( 36,8)),
			1863 => std_logic_vector(to_unsigned( 214,8)),
			1864 => std_logic_vector(to_unsigned( 131,8)),
			1865 => std_logic_vector(to_unsigned( 40,8)),
			1866 => std_logic_vector(to_unsigned( 58,8)),
			1867 => std_logic_vector(to_unsigned( 2,8)),
			1868 => std_logic_vector(to_unsigned( 250,8)),
			1869 => std_logic_vector(to_unsigned( 60,8)),
			1870 => std_logic_vector(to_unsigned( 234,8)),
			1871 => std_logic_vector(to_unsigned( 67,8)),
			1872 => std_logic_vector(to_unsigned( 70,8)),
			1873 => std_logic_vector(to_unsigned( 16,8)),
			1874 => std_logic_vector(to_unsigned( 12,8)),
			1875 => std_logic_vector(to_unsigned( 233,8)),
			1876 => std_logic_vector(to_unsigned( 112,8)),
			1877 => std_logic_vector(to_unsigned( 253,8)),
			1878 => std_logic_vector(to_unsigned( 251,8)),
			1879 => std_logic_vector(to_unsigned( 16,8)),
			1880 => std_logic_vector(to_unsigned( 126,8)),
			1881 => std_logic_vector(to_unsigned( 242,8)),
			1882 => std_logic_vector(to_unsigned( 146,8)),
			1883 => std_logic_vector(to_unsigned( 156,8)),
			1884 => std_logic_vector(to_unsigned( 160,8)),
			1885 => std_logic_vector(to_unsigned( 218,8)),
			1886 => std_logic_vector(to_unsigned( 138,8)),
			1887 => std_logic_vector(to_unsigned( 149,8)),
			1888 => std_logic_vector(to_unsigned( 140,8)),
			1889 => std_logic_vector(to_unsigned( 126,8)),
			1890 => std_logic_vector(to_unsigned( 224,8)),
			1891 => std_logic_vector(to_unsigned( 135,8)),
			1892 => std_logic_vector(to_unsigned( 238,8)),
			1893 => std_logic_vector(to_unsigned( 124,8)),
			1894 => std_logic_vector(to_unsigned( 54,8)),
			1895 => std_logic_vector(to_unsigned( 113,8)),
			1896 => std_logic_vector(to_unsigned( 106,8)),
			1897 => std_logic_vector(to_unsigned( 236,8)),
			1898 => std_logic_vector(to_unsigned( 46,8)),
			1899 => std_logic_vector(to_unsigned( 85,8)),
			1900 => std_logic_vector(to_unsigned( 170,8)),
			1901 => std_logic_vector(to_unsigned( 6,8)),
			1902 => std_logic_vector(to_unsigned( 194,8)),
			1903 => std_logic_vector(to_unsigned( 18,8)),
			1904 => std_logic_vector(to_unsigned( 234,8)),
			1905 => std_logic_vector(to_unsigned( 17,8)),
			1906 => std_logic_vector(to_unsigned( 20,8)),
			1907 => std_logic_vector(to_unsigned( 160,8)),
			1908 => std_logic_vector(to_unsigned( 202,8)),
			1909 => std_logic_vector(to_unsigned( 170,8)),
			1910 => std_logic_vector(to_unsigned( 88,8)),
			1911 => std_logic_vector(to_unsigned( 205,8)),
			1912 => std_logic_vector(to_unsigned( 219,8)),
			1913 => std_logic_vector(to_unsigned( 176,8)),
			1914 => std_logic_vector(to_unsigned( 67,8)),
			1915 => std_logic_vector(to_unsigned( 180,8)),
			1916 => std_logic_vector(to_unsigned( 236,8)),
			1917 => std_logic_vector(to_unsigned( 172,8)),
			1918 => std_logic_vector(to_unsigned( 13,8)),
			1919 => std_logic_vector(to_unsigned( 215,8)),
			1920 => std_logic_vector(to_unsigned( 23,8)),
			1921 => std_logic_vector(to_unsigned( 241,8)),
			1922 => std_logic_vector(to_unsigned( 62,8)),
			1923 => std_logic_vector(to_unsigned( 68,8)),
			1924 => std_logic_vector(to_unsigned( 172,8)),
			1925 => std_logic_vector(to_unsigned( 13,8)),
			1926 => std_logic_vector(to_unsigned( 249,8)),
			1927 => std_logic_vector(to_unsigned( 21,8)),
			1928 => std_logic_vector(to_unsigned( 106,8)),
			1929 => std_logic_vector(to_unsigned( 211,8)),
			1930 => std_logic_vector(to_unsigned( 41,8)),
			1931 => std_logic_vector(to_unsigned( 52,8)),
			1932 => std_logic_vector(to_unsigned( 121,8)),
			1933 => std_logic_vector(to_unsigned( 120,8)),
			1934 => std_logic_vector(to_unsigned( 36,8)),
			1935 => std_logic_vector(to_unsigned( 146,8)),
			1936 => std_logic_vector(to_unsigned( 245,8)),
			1937 => std_logic_vector(to_unsigned( 108,8)),
			1938 => std_logic_vector(to_unsigned( 68,8)),
			1939 => std_logic_vector(to_unsigned( 141,8)),
			1940 => std_logic_vector(to_unsigned( 18,8)),
			1941 => std_logic_vector(to_unsigned( 74,8)),
			1942 => std_logic_vector(to_unsigned( 220,8)),
			1943 => std_logic_vector(to_unsigned( 224,8)),
			1944 => std_logic_vector(to_unsigned( 14,8)),
			1945 => std_logic_vector(to_unsigned( 249,8)),
			1946 => std_logic_vector(to_unsigned( 190,8)),
			1947 => std_logic_vector(to_unsigned( 59,8)),
			1948 => std_logic_vector(to_unsigned( 196,8)),
			1949 => std_logic_vector(to_unsigned( 255,8)),
			1950 => std_logic_vector(to_unsigned( 33,8)),
			1951 => std_logic_vector(to_unsigned( 52,8)),
			1952 => std_logic_vector(to_unsigned( 79,8)),
			1953 => std_logic_vector(to_unsigned( 232,8)),
			1954 => std_logic_vector(to_unsigned( 130,8)),
			1955 => std_logic_vector(to_unsigned( 107,8)),
			1956 => std_logic_vector(to_unsigned( 230,8)),
			1957 => std_logic_vector(to_unsigned( 41,8)),
			1958 => std_logic_vector(to_unsigned( 157,8)),
			1959 => std_logic_vector(to_unsigned( 145,8)),
			1960 => std_logic_vector(to_unsigned( 114,8)),
			1961 => std_logic_vector(to_unsigned( 151,8)),
			1962 => std_logic_vector(to_unsigned( 137,8)),
			1963 => std_logic_vector(to_unsigned( 240,8)),
			1964 => std_logic_vector(to_unsigned( 141,8)),
			1965 => std_logic_vector(to_unsigned( 229,8)),
			1966 => std_logic_vector(to_unsigned( 94,8)),
			1967 => std_logic_vector(to_unsigned( 167,8)),
			1968 => std_logic_vector(to_unsigned( 208,8)),
			1969 => std_logic_vector(to_unsigned( 152,8)),
			1970 => std_logic_vector(to_unsigned( 12,8)),
			1971 => std_logic_vector(to_unsigned( 232,8)),
			1972 => std_logic_vector(to_unsigned( 123,8)),
			1973 => std_logic_vector(to_unsigned( 133,8)),
			1974 => std_logic_vector(to_unsigned( 181,8)),
			1975 => std_logic_vector(to_unsigned( 21,8)),
			1976 => std_logic_vector(to_unsigned( 159,8)),
			1977 => std_logic_vector(to_unsigned( 175,8)),
			1978 => std_logic_vector(to_unsigned( 108,8)),
			1979 => std_logic_vector(to_unsigned( 82,8)),
			1980 => std_logic_vector(to_unsigned( 103,8)),
			1981 => std_logic_vector(to_unsigned( 23,8)),
			1982 => std_logic_vector(to_unsigned( 219,8)),
			1983 => std_logic_vector(to_unsigned( 68,8)),
			1984 => std_logic_vector(to_unsigned( 51,8)),
			1985 => std_logic_vector(to_unsigned( 248,8)),
			1986 => std_logic_vector(to_unsigned( 172,8)),
			1987 => std_logic_vector(to_unsigned( 204,8)),
			1988 => std_logic_vector(to_unsigned( 21,8)),
			1989 => std_logic_vector(to_unsigned( 240,8)),
			1990 => std_logic_vector(to_unsigned( 165,8)),
			1991 => std_logic_vector(to_unsigned( 47,8)),
			1992 => std_logic_vector(to_unsigned( 117,8)),
			1993 => std_logic_vector(to_unsigned( 54,8)),
			1994 => std_logic_vector(to_unsigned( 232,8)),
			1995 => std_logic_vector(to_unsigned( 105,8)),
			1996 => std_logic_vector(to_unsigned( 231,8)),
			1997 => std_logic_vector(to_unsigned( 174,8)),
			1998 => std_logic_vector(to_unsigned( 41,8)),
			1999 => std_logic_vector(to_unsigned( 224,8)),
			2000 => std_logic_vector(to_unsigned( 82,8)),
			2001 => std_logic_vector(to_unsigned( 234,8)),
			2002 => std_logic_vector(to_unsigned( 65,8)),
			2003 => std_logic_vector(to_unsigned( 223,8)),
			2004 => std_logic_vector(to_unsigned( 156,8)),
			2005 => std_logic_vector(to_unsigned( 14,8)),
			2006 => std_logic_vector(to_unsigned( 217,8)),
			2007 => std_logic_vector(to_unsigned( 127,8)),
			2008 => std_logic_vector(to_unsigned( 41,8)),
			2009 => std_logic_vector(to_unsigned( 122,8)),
			2010 => std_logic_vector(to_unsigned( 94,8)),
			2011 => std_logic_vector(to_unsigned( 243,8)),
			2012 => std_logic_vector(to_unsigned( 145,8)),
			2013 => std_logic_vector(to_unsigned( 203,8)),
			2014 => std_logic_vector(to_unsigned( 49,8)),
			2015 => std_logic_vector(to_unsigned( 126,8)),
			2016 => std_logic_vector(to_unsigned( 30,8)),
			2017 => std_logic_vector(to_unsigned( 82,8)),
			2018 => std_logic_vector(to_unsigned( 252,8)),
			2019 => std_logic_vector(to_unsigned( 4,8)),
			2020 => std_logic_vector(to_unsigned( 131,8)),
			2021 => std_logic_vector(to_unsigned( 144,8)),
			2022 => std_logic_vector(to_unsigned( 25,8)),
			2023 => std_logic_vector(to_unsigned( 32,8)),
			2024 => std_logic_vector(to_unsigned( 140,8)),
			2025 => std_logic_vector(to_unsigned( 120,8)),
			2026 => std_logic_vector(to_unsigned( 237,8)),
			2027 => std_logic_vector(to_unsigned( 56,8)),
			2028 => std_logic_vector(to_unsigned( 189,8)),
			2029 => std_logic_vector(to_unsigned( 198,8)),
			2030 => std_logic_vector(to_unsigned( 166,8)),
			2031 => std_logic_vector(to_unsigned( 144,8)),
			2032 => std_logic_vector(to_unsigned( 218,8)),
			2033 => std_logic_vector(to_unsigned( 91,8)),
			2034 => std_logic_vector(to_unsigned( 193,8)),
			2035 => std_logic_vector(to_unsigned( 225,8)),
			2036 => std_logic_vector(to_unsigned( 40,8)),
			2037 => std_logic_vector(to_unsigned( 252,8)),
			2038 => std_logic_vector(to_unsigned( 123,8)),
			2039 => std_logic_vector(to_unsigned( 223,8)),
			2040 => std_logic_vector(to_unsigned( 9,8)),
			2041 => std_logic_vector(to_unsigned( 113,8)),
			2042 => std_logic_vector(to_unsigned( 4,8)),
			2043 => std_logic_vector(to_unsigned( 107,8)),
			2044 => std_logic_vector(to_unsigned( 145,8)),
			2045 => std_logic_vector(to_unsigned( 217,8)),
			2046 => std_logic_vector(to_unsigned( 250,8)),
			2047 => std_logic_vector(to_unsigned( 253,8)),
			2048 => std_logic_vector(to_unsigned( 195,8)),
			2049 => std_logic_vector(to_unsigned( 109,8)),
			2050 => std_logic_vector(to_unsigned( 190,8)),
			2051 => std_logic_vector(to_unsigned( 95,8)),
			2052 => std_logic_vector(to_unsigned( 254,8)),
			2053 => std_logic_vector(to_unsigned( 233,8)),
			2054 => std_logic_vector(to_unsigned( 215,8)),
			2055 => std_logic_vector(to_unsigned( 11,8)),
			2056 => std_logic_vector(to_unsigned( 83,8)),
			2057 => std_logic_vector(to_unsigned( 81,8)),
			2058 => std_logic_vector(to_unsigned( 24,8)),
			2059 => std_logic_vector(to_unsigned( 156,8)),
			2060 => std_logic_vector(to_unsigned( 197,8)),
			2061 => std_logic_vector(to_unsigned( 239,8)),
			2062 => std_logic_vector(to_unsigned( 88,8)),
			2063 => std_logic_vector(to_unsigned( 204,8)),
			2064 => std_logic_vector(to_unsigned( 140,8)),
			2065 => std_logic_vector(to_unsigned( 161,8)),
			2066 => std_logic_vector(to_unsigned( 122,8)),
			2067 => std_logic_vector(to_unsigned( 41,8)),
			2068 => std_logic_vector(to_unsigned( 89,8)),
			2069 => std_logic_vector(to_unsigned( 202,8)),
			2070 => std_logic_vector(to_unsigned( 217,8)),
			2071 => std_logic_vector(to_unsigned( 94,8)),
			2072 => std_logic_vector(to_unsigned( 170,8)),
			2073 => std_logic_vector(to_unsigned( 9,8)),
			2074 => std_logic_vector(to_unsigned( 232,8)),
			2075 => std_logic_vector(to_unsigned( 41,8)),
			2076 => std_logic_vector(to_unsigned( 29,8)),
			2077 => std_logic_vector(to_unsigned( 71,8)),
			2078 => std_logic_vector(to_unsigned( 187,8)),
			2079 => std_logic_vector(to_unsigned( 161,8)),
			2080 => std_logic_vector(to_unsigned( 108,8)),
			2081 => std_logic_vector(to_unsigned( 178,8)),
			2082 => std_logic_vector(to_unsigned( 225,8)),
			2083 => std_logic_vector(to_unsigned( 248,8)),
			2084 => std_logic_vector(to_unsigned( 18,8)),
			2085 => std_logic_vector(to_unsigned( 240,8)),
			2086 => std_logic_vector(to_unsigned( 133,8)),
			2087 => std_logic_vector(to_unsigned( 96,8)),
			2088 => std_logic_vector(to_unsigned( 78,8)),
			2089 => std_logic_vector(to_unsigned( 204,8)),
			2090 => std_logic_vector(to_unsigned( 31,8)),
			2091 => std_logic_vector(to_unsigned( 145,8)),
			2092 => std_logic_vector(to_unsigned( 218,8)),
			2093 => std_logic_vector(to_unsigned( 67,8)),
			2094 => std_logic_vector(to_unsigned( 30,8)),
			2095 => std_logic_vector(to_unsigned( 182,8)),
			2096 => std_logic_vector(to_unsigned( 134,8)),
			2097 => std_logic_vector(to_unsigned( 29,8)),
			2098 => std_logic_vector(to_unsigned( 121,8)),
			2099 => std_logic_vector(to_unsigned( 98,8)),
			2100 => std_logic_vector(to_unsigned( 28,8)),
			2101 => std_logic_vector(to_unsigned( 191,8)),
			2102 => std_logic_vector(to_unsigned( 240,8)),
			2103 => std_logic_vector(to_unsigned( 214,8)),
			2104 => std_logic_vector(to_unsigned( 55,8)),
			2105 => std_logic_vector(to_unsigned( 210,8)),
			2106 => std_logic_vector(to_unsigned( 122,8)),
			2107 => std_logic_vector(to_unsigned( 50,8)),
			2108 => std_logic_vector(to_unsigned( 216,8)),
			2109 => std_logic_vector(to_unsigned( 38,8)),
			2110 => std_logic_vector(to_unsigned( 225,8)),
			2111 => std_logic_vector(to_unsigned( 95,8)),
			2112 => std_logic_vector(to_unsigned( 11,8)),
			2113 => std_logic_vector(to_unsigned( 219,8)),
			2114 => std_logic_vector(to_unsigned( 254,8)),
			2115 => std_logic_vector(to_unsigned( 167,8)),
			2116 => std_logic_vector(to_unsigned( 248,8)),
			2117 => std_logic_vector(to_unsigned( 238,8)),
			2118 => std_logic_vector(to_unsigned( 107,8)),
			2119 => std_logic_vector(to_unsigned( 1,8)),
			2120 => std_logic_vector(to_unsigned( 187,8)),
			2121 => std_logic_vector(to_unsigned( 20,8)),
			2122 => std_logic_vector(to_unsigned( 13,8)),
			2123 => std_logic_vector(to_unsigned( 151,8)),
			2124 => std_logic_vector(to_unsigned( 159,8)),
			2125 => std_logic_vector(to_unsigned( 101,8)),
			2126 => std_logic_vector(to_unsigned( 169,8)),
			2127 => std_logic_vector(to_unsigned( 203,8)),
			2128 => std_logic_vector(to_unsigned( 85,8)),
			2129 => std_logic_vector(to_unsigned( 17,8)),
			2130 => std_logic_vector(to_unsigned( 194,8)),
			2131 => std_logic_vector(to_unsigned( 11,8)),
			2132 => std_logic_vector(to_unsigned( 177,8)),
			2133 => std_logic_vector(to_unsigned( 246,8)),
			2134 => std_logic_vector(to_unsigned( 152,8)),
			2135 => std_logic_vector(to_unsigned( 183,8)),
			2136 => std_logic_vector(to_unsigned( 3,8)),
			2137 => std_logic_vector(to_unsigned( 99,8)),
			2138 => std_logic_vector(to_unsigned( 63,8)),
			2139 => std_logic_vector(to_unsigned( 123,8)),
			2140 => std_logic_vector(to_unsigned( 104,8)),
			2141 => std_logic_vector(to_unsigned( 39,8)),
			2142 => std_logic_vector(to_unsigned( 88,8)),
			2143 => std_logic_vector(to_unsigned( 37,8)),
			2144 => std_logic_vector(to_unsigned( 118,8)),
			2145 => std_logic_vector(to_unsigned( 99,8)),
			2146 => std_logic_vector(to_unsigned( 87,8)),
			2147 => std_logic_vector(to_unsigned( 34,8)),
			2148 => std_logic_vector(to_unsigned( 68,8)),
			2149 => std_logic_vector(to_unsigned( 75,8)),
			2150 => std_logic_vector(to_unsigned( 18,8)),
			2151 => std_logic_vector(to_unsigned( 92,8)),
			2152 => std_logic_vector(to_unsigned( 111,8)),
			2153 => std_logic_vector(to_unsigned( 208,8)),
			2154 => std_logic_vector(to_unsigned( 53,8)),
			2155 => std_logic_vector(to_unsigned( 43,8)),
			2156 => std_logic_vector(to_unsigned( 192,8)),
			2157 => std_logic_vector(to_unsigned( 217,8)),
			2158 => std_logic_vector(to_unsigned( 12,8)),
			2159 => std_logic_vector(to_unsigned( 39,8)),
			2160 => std_logic_vector(to_unsigned( 86,8)),
			2161 => std_logic_vector(to_unsigned( 144,8)),
			2162 => std_logic_vector(to_unsigned( 177,8)),
			2163 => std_logic_vector(to_unsigned( 162,8)),
			2164 => std_logic_vector(to_unsigned( 41,8)),
			2165 => std_logic_vector(to_unsigned( 198,8)),
			2166 => std_logic_vector(to_unsigned( 11,8)),
			2167 => std_logic_vector(to_unsigned( 18,8)),
			2168 => std_logic_vector(to_unsigned( 93,8)),
			2169 => std_logic_vector(to_unsigned( 211,8)),
			2170 => std_logic_vector(to_unsigned( 111,8)),
			2171 => std_logic_vector(to_unsigned( 145,8)),
			2172 => std_logic_vector(to_unsigned( 16,8)),
			2173 => std_logic_vector(to_unsigned( 200,8)),
			2174 => std_logic_vector(to_unsigned( 41,8)),
			2175 => std_logic_vector(to_unsigned( 219,8)),
			2176 => std_logic_vector(to_unsigned( 139,8)),
			2177 => std_logic_vector(to_unsigned( 150,8)),
			2178 => std_logic_vector(to_unsigned( 238,8)),
			2179 => std_logic_vector(to_unsigned( 164,8)),
			2180 => std_logic_vector(to_unsigned( 156,8)),
			2181 => std_logic_vector(to_unsigned( 77,8)),
			2182 => std_logic_vector(to_unsigned( 202,8)),
			2183 => std_logic_vector(to_unsigned( 150,8)),
			2184 => std_logic_vector(to_unsigned( 113,8)),
			2185 => std_logic_vector(to_unsigned( 135,8)),
			2186 => std_logic_vector(to_unsigned( 137,8)),
			2187 => std_logic_vector(to_unsigned( 241,8)),
			2188 => std_logic_vector(to_unsigned( 3,8)),
			2189 => std_logic_vector(to_unsigned( 146,8)),
			2190 => std_logic_vector(to_unsigned( 190,8)),
			2191 => std_logic_vector(to_unsigned( 43,8)),
			2192 => std_logic_vector(to_unsigned( 203,8)),
			2193 => std_logic_vector(to_unsigned( 205,8)),
			2194 => std_logic_vector(to_unsigned( 252,8)),
			2195 => std_logic_vector(to_unsigned( 103,8)),
			2196 => std_logic_vector(to_unsigned( 170,8)),
			2197 => std_logic_vector(to_unsigned( 167,8)),
			2198 => std_logic_vector(to_unsigned( 164,8)),
			2199 => std_logic_vector(to_unsigned( 10,8)),
			2200 => std_logic_vector(to_unsigned( 85,8)),
			2201 => std_logic_vector(to_unsigned( 58,8)),
			2202 => std_logic_vector(to_unsigned( 108,8)),
			2203 => std_logic_vector(to_unsigned( 4,8)),
			2204 => std_logic_vector(to_unsigned( 221,8)),
			2205 => std_logic_vector(to_unsigned( 225,8)),
			2206 => std_logic_vector(to_unsigned( 161,8)),
			2207 => std_logic_vector(to_unsigned( 31,8)),
			2208 => std_logic_vector(to_unsigned( 18,8)),
			2209 => std_logic_vector(to_unsigned( 110,8)),
			2210 => std_logic_vector(to_unsigned( 222,8)),
			2211 => std_logic_vector(to_unsigned( 20,8)),
			2212 => std_logic_vector(to_unsigned( 11,8)),
			2213 => std_logic_vector(to_unsigned( 110,8)),
			2214 => std_logic_vector(to_unsigned( 147,8)),
			2215 => std_logic_vector(to_unsigned( 137,8)),
			2216 => std_logic_vector(to_unsigned( 174,8)),
			2217 => std_logic_vector(to_unsigned( 3,8)),
			2218 => std_logic_vector(to_unsigned( 17,8)),
			2219 => std_logic_vector(to_unsigned( 151,8)),
			2220 => std_logic_vector(to_unsigned( 71,8)),
			2221 => std_logic_vector(to_unsigned( 234,8)),
			2222 => std_logic_vector(to_unsigned( 54,8)),
			2223 => std_logic_vector(to_unsigned( 115,8)),
			2224 => std_logic_vector(to_unsigned( 97,8)),
			2225 => std_logic_vector(to_unsigned( 235,8)),
			2226 => std_logic_vector(to_unsigned( 59,8)),
			2227 => std_logic_vector(to_unsigned( 21,8)),
			2228 => std_logic_vector(to_unsigned( 87,8)),
			2229 => std_logic_vector(to_unsigned( 248,8)),
			2230 => std_logic_vector(to_unsigned( 201,8)),
			2231 => std_logic_vector(to_unsigned( 62,8)),
			2232 => std_logic_vector(to_unsigned( 68,8)),
			2233 => std_logic_vector(to_unsigned( 187,8)),
			2234 => std_logic_vector(to_unsigned( 12,8)),
			2235 => std_logic_vector(to_unsigned( 49,8)),
			2236 => std_logic_vector(to_unsigned( 115,8)),
			2237 => std_logic_vector(to_unsigned( 167,8)),
			2238 => std_logic_vector(to_unsigned( 19,8)),
			2239 => std_logic_vector(to_unsigned( 108,8)),
			2240 => std_logic_vector(to_unsigned( 239,8)),
			2241 => std_logic_vector(to_unsigned( 225,8)),
			2242 => std_logic_vector(to_unsigned( 252,8)),
			2243 => std_logic_vector(to_unsigned( 217,8)),
			2244 => std_logic_vector(to_unsigned( 198,8)),
			2245 => std_logic_vector(to_unsigned( 10,8)),
			2246 => std_logic_vector(to_unsigned( 236,8)),
			2247 => std_logic_vector(to_unsigned( 55,8)),
			2248 => std_logic_vector(to_unsigned( 91,8)),
			2249 => std_logic_vector(to_unsigned( 83,8)),
			2250 => std_logic_vector(to_unsigned( 90,8)),
			2251 => std_logic_vector(to_unsigned( 87,8)),
			2252 => std_logic_vector(to_unsigned( 236,8)),
			2253 => std_logic_vector(to_unsigned( 23,8)),
			2254 => std_logic_vector(to_unsigned( 170,8)),
			2255 => std_logic_vector(to_unsigned( 184,8)),
			2256 => std_logic_vector(to_unsigned( 121,8)),
			2257 => std_logic_vector(to_unsigned( 25,8)),
			2258 => std_logic_vector(to_unsigned( 94,8)),
			2259 => std_logic_vector(to_unsigned( 90,8)),
			2260 => std_logic_vector(to_unsigned( 215,8)),
			2261 => std_logic_vector(to_unsigned( 4,8)),
			2262 => std_logic_vector(to_unsigned( 136,8)),
			2263 => std_logic_vector(to_unsigned( 126,8)),
			2264 => std_logic_vector(to_unsigned( 109,8)),
			2265 => std_logic_vector(to_unsigned( 55,8)),
			2266 => std_logic_vector(to_unsigned( 116,8)),
			2267 => std_logic_vector(to_unsigned( 58,8)),
			2268 => std_logic_vector(to_unsigned( 114,8)),
			2269 => std_logic_vector(to_unsigned( 149,8)),
			2270 => std_logic_vector(to_unsigned( 61,8)),
			2271 => std_logic_vector(to_unsigned( 52,8)),
			2272 => std_logic_vector(to_unsigned( 65,8)),
			2273 => std_logic_vector(to_unsigned( 157,8)),
			2274 => std_logic_vector(to_unsigned( 43,8)),
			2275 => std_logic_vector(to_unsigned( 229,8)),
			2276 => std_logic_vector(to_unsigned( 195,8)),
			2277 => std_logic_vector(to_unsigned( 44,8)),
			2278 => std_logic_vector(to_unsigned( 221,8)),
			2279 => std_logic_vector(to_unsigned( 59,8)),
			2280 => std_logic_vector(to_unsigned( 78,8)),
			2281 => std_logic_vector(to_unsigned( 13,8)),
			2282 => std_logic_vector(to_unsigned( 74,8)),
			2283 => std_logic_vector(to_unsigned( 209,8)),
			2284 => std_logic_vector(to_unsigned( 106,8)),
			2285 => std_logic_vector(to_unsigned( 135,8)),
			2286 => std_logic_vector(to_unsigned( 142,8)),
			2287 => std_logic_vector(to_unsigned( 223,8)),
			2288 => std_logic_vector(to_unsigned( 12,8)),
			2289 => std_logic_vector(to_unsigned( 20,8)),
			2290 => std_logic_vector(to_unsigned( 83,8)),
			2291 => std_logic_vector(to_unsigned( 193,8)),
			2292 => std_logic_vector(to_unsigned( 44,8)),
			2293 => std_logic_vector(to_unsigned( 8,8)),
			2294 => std_logic_vector(to_unsigned( 246,8)),
			2295 => std_logic_vector(to_unsigned( 141,8)),
			2296 => std_logic_vector(to_unsigned( 168,8)),
			2297 => std_logic_vector(to_unsigned( 25,8)),
			2298 => std_logic_vector(to_unsigned( 189,8)),
			2299 => std_logic_vector(to_unsigned( 105,8)),
			2300 => std_logic_vector(to_unsigned( 33,8)),
			2301 => std_logic_vector(to_unsigned( 88,8)),
			2302 => std_logic_vector(to_unsigned( 153,8)),
			2303 => std_logic_vector(to_unsigned( 145,8)),
			2304 => std_logic_vector(to_unsigned( 157,8)),
			2305 => std_logic_vector(to_unsigned( 220,8)),
			2306 => std_logic_vector(to_unsigned( 2,8)),
			2307 => std_logic_vector(to_unsigned( 17,8)),
			2308 => std_logic_vector(to_unsigned( 81,8)),
			2309 => std_logic_vector(to_unsigned( 178,8)),
			2310 => std_logic_vector(to_unsigned( 205,8)),
			2311 => std_logic_vector(to_unsigned( 20,8)),
			2312 => std_logic_vector(to_unsigned( 55,8)),
			2313 => std_logic_vector(to_unsigned( 244,8)),
			2314 => std_logic_vector(to_unsigned( 191,8)),
			2315 => std_logic_vector(to_unsigned( 129,8)),
			2316 => std_logic_vector(to_unsigned( 242,8)),
			2317 => std_logic_vector(to_unsigned( 245,8)),
			2318 => std_logic_vector(to_unsigned( 181,8)),
			2319 => std_logic_vector(to_unsigned( 204,8)),
			2320 => std_logic_vector(to_unsigned( 85,8)),
			2321 => std_logic_vector(to_unsigned( 171,8)),
			2322 => std_logic_vector(to_unsigned( 108,8)),
			2323 => std_logic_vector(to_unsigned( 9,8)),
			2324 => std_logic_vector(to_unsigned( 11,8)),
			2325 => std_logic_vector(to_unsigned( 193,8)),
			2326 => std_logic_vector(to_unsigned( 5,8)),
			2327 => std_logic_vector(to_unsigned( 234,8)),
			2328 => std_logic_vector(to_unsigned( 221,8)),
			2329 => std_logic_vector(to_unsigned( 5,8)),
			2330 => std_logic_vector(to_unsigned( 187,8)),
			2331 => std_logic_vector(to_unsigned( 168,8)),
			2332 => std_logic_vector(to_unsigned( 64,8)),
			2333 => std_logic_vector(to_unsigned( 126,8)),
			2334 => std_logic_vector(to_unsigned( 6,8)),
			2335 => std_logic_vector(to_unsigned( 151,8)),
			2336 => std_logic_vector(to_unsigned( 71,8)),
			2337 => std_logic_vector(to_unsigned( 182,8)),
			2338 => std_logic_vector(to_unsigned( 65,8)),
			2339 => std_logic_vector(to_unsigned( 90,8)),
			2340 => std_logic_vector(to_unsigned( 108,8)),
			2341 => std_logic_vector(to_unsigned( 148,8)),
			2342 => std_logic_vector(to_unsigned( 75,8)),
			2343 => std_logic_vector(to_unsigned( 220,8)),
			2344 => std_logic_vector(to_unsigned( 158,8)),
			2345 => std_logic_vector(to_unsigned( 52,8)),
			2346 => std_logic_vector(to_unsigned( 205,8)),
			2347 => std_logic_vector(to_unsigned( 2,8)),
			2348 => std_logic_vector(to_unsigned( 141,8)),
			2349 => std_logic_vector(to_unsigned( 124,8)),
			2350 => std_logic_vector(to_unsigned( 61,8)),
			2351 => std_logic_vector(to_unsigned( 173,8)),
			2352 => std_logic_vector(to_unsigned( 245,8)),
			2353 => std_logic_vector(to_unsigned( 119,8)),
			2354 => std_logic_vector(to_unsigned( 91,8)),
			2355 => std_logic_vector(to_unsigned( 33,8)),
			2356 => std_logic_vector(to_unsigned( 22,8)),
			2357 => std_logic_vector(to_unsigned( 244,8)),
			2358 => std_logic_vector(to_unsigned( 226,8)),
			2359 => std_logic_vector(to_unsigned( 175,8)),
			2360 => std_logic_vector(to_unsigned( 151,8)),
			2361 => std_logic_vector(to_unsigned( 241,8)),
			2362 => std_logic_vector(to_unsigned( 197,8)),
			2363 => std_logic_vector(to_unsigned( 7,8)),
			2364 => std_logic_vector(to_unsigned( 95,8)),
			2365 => std_logic_vector(to_unsigned( 215,8)),
			2366 => std_logic_vector(to_unsigned( 150,8)),
			2367 => std_logic_vector(to_unsigned( 247,8)),
			2368 => std_logic_vector(to_unsigned( 92,8)),
			2369 => std_logic_vector(to_unsigned( 3,8)),
			2370 => std_logic_vector(to_unsigned( 156,8)),
			2371 => std_logic_vector(to_unsigned( 49,8)),
			2372 => std_logic_vector(to_unsigned( 119,8)),
			2373 => std_logic_vector(to_unsigned( 132,8)),
			2374 => std_logic_vector(to_unsigned( 254,8)),
			2375 => std_logic_vector(to_unsigned( 244,8)),
			2376 => std_logic_vector(to_unsigned( 199,8)),
			2377 => std_logic_vector(to_unsigned( 3,8)),
			2378 => std_logic_vector(to_unsigned( 163,8)),
			2379 => std_logic_vector(to_unsigned( 175,8)),
			2380 => std_logic_vector(to_unsigned( 217,8)),
			2381 => std_logic_vector(to_unsigned( 29,8)),
			2382 => std_logic_vector(to_unsigned( 143,8)),
			2383 => std_logic_vector(to_unsigned( 142,8)),
			2384 => std_logic_vector(to_unsigned( 11,8)),
			2385 => std_logic_vector(to_unsigned( 79,8)),
			2386 => std_logic_vector(to_unsigned( 123,8)),
			2387 => std_logic_vector(to_unsigned( 182,8)),
			2388 => std_logic_vector(to_unsigned( 33,8)),
			2389 => std_logic_vector(to_unsigned( 43,8)),
			2390 => std_logic_vector(to_unsigned( 14,8)),
			2391 => std_logic_vector(to_unsigned( 185,8)),
			2392 => std_logic_vector(to_unsigned( 138,8)),
			2393 => std_logic_vector(to_unsigned( 68,8)),
			2394 => std_logic_vector(to_unsigned( 19,8)),
			2395 => std_logic_vector(to_unsigned( 113,8)),
			2396 => std_logic_vector(to_unsigned( 76,8)),
			2397 => std_logic_vector(to_unsigned( 114,8)),
			2398 => std_logic_vector(to_unsigned( 140,8)),
			2399 => std_logic_vector(to_unsigned( 203,8)),
			2400 => std_logic_vector(to_unsigned( 196,8)),
			2401 => std_logic_vector(to_unsigned( 176,8)),
			2402 => std_logic_vector(to_unsigned( 232,8)),
			2403 => std_logic_vector(to_unsigned( 12,8)),
			2404 => std_logic_vector(to_unsigned( 245,8)),
			2405 => std_logic_vector(to_unsigned( 135,8)),
			2406 => std_logic_vector(to_unsigned( 22,8)),
			2407 => std_logic_vector(to_unsigned( 209,8)),
			2408 => std_logic_vector(to_unsigned( 115,8)),
			2409 => std_logic_vector(to_unsigned( 82,8)),
			2410 => std_logic_vector(to_unsigned( 58,8)),
			2411 => std_logic_vector(to_unsigned( 114,8)),
			2412 => std_logic_vector(to_unsigned( 233,8)),
			2413 => std_logic_vector(to_unsigned( 203,8)),
			2414 => std_logic_vector(to_unsigned( 197,8)),
			2415 => std_logic_vector(to_unsigned( 26,8)),
			2416 => std_logic_vector(to_unsigned( 185,8)),
			2417 => std_logic_vector(to_unsigned( 110,8)),
			2418 => std_logic_vector(to_unsigned( 97,8)),
			2419 => std_logic_vector(to_unsigned( 96,8)),
			2420 => std_logic_vector(to_unsigned( 162,8)),
			2421 => std_logic_vector(to_unsigned( 171,8)),
			2422 => std_logic_vector(to_unsigned( 104,8)),
			2423 => std_logic_vector(to_unsigned( 79,8)),
			2424 => std_logic_vector(to_unsigned( 18,8)),
			2425 => std_logic_vector(to_unsigned( 218,8)),
			2426 => std_logic_vector(to_unsigned( 48,8)),
			2427 => std_logic_vector(to_unsigned( 7,8)),
			2428 => std_logic_vector(to_unsigned( 120,8)),
			2429 => std_logic_vector(to_unsigned( 228,8)),
			2430 => std_logic_vector(to_unsigned( 82,8)),
			2431 => std_logic_vector(to_unsigned( 104,8)),
			2432 => std_logic_vector(to_unsigned( 30,8)),
			2433 => std_logic_vector(to_unsigned( 45,8)),
			2434 => std_logic_vector(to_unsigned( 11,8)),
			2435 => std_logic_vector(to_unsigned( 120,8)),
			2436 => std_logic_vector(to_unsigned( 16,8)),
			2437 => std_logic_vector(to_unsigned( 129,8)),
			2438 => std_logic_vector(to_unsigned( 235,8)),
			2439 => std_logic_vector(to_unsigned( 191,8)),
			2440 => std_logic_vector(to_unsigned( 107,8)),
			2441 => std_logic_vector(to_unsigned( 4,8)),
			2442 => std_logic_vector(to_unsigned( 147,8)),
			2443 => std_logic_vector(to_unsigned( 252,8)),
			2444 => std_logic_vector(to_unsigned( 146,8)),
			2445 => std_logic_vector(to_unsigned( 126,8)),
			2446 => std_logic_vector(to_unsigned( 31,8)),
			2447 => std_logic_vector(to_unsigned( 18,8)),
			2448 => std_logic_vector(to_unsigned( 219,8)),
			2449 => std_logic_vector(to_unsigned( 42,8)),
			2450 => std_logic_vector(to_unsigned( 195,8)),
			2451 => std_logic_vector(to_unsigned( 192,8)),
			2452 => std_logic_vector(to_unsigned( 187,8)),
			2453 => std_logic_vector(to_unsigned( 235,8)),
			2454 => std_logic_vector(to_unsigned( 117,8)),
			2455 => std_logic_vector(to_unsigned( 61,8)),
			2456 => std_logic_vector(to_unsigned( 59,8)),
			2457 => std_logic_vector(to_unsigned( 37,8)),
			2458 => std_logic_vector(to_unsigned( 32,8)),
			2459 => std_logic_vector(to_unsigned( 139,8)),
			2460 => std_logic_vector(to_unsigned( 23,8)),
			2461 => std_logic_vector(to_unsigned( 9,8)),
			2462 => std_logic_vector(to_unsigned( 191,8)),
			2463 => std_logic_vector(to_unsigned( 55,8)),
			2464 => std_logic_vector(to_unsigned( 113,8)),
			2465 => std_logic_vector(to_unsigned( 180,8)),
			2466 => std_logic_vector(to_unsigned( 168,8)),
			2467 => std_logic_vector(to_unsigned( 124,8)),
			2468 => std_logic_vector(to_unsigned( 105,8)),
			2469 => std_logic_vector(to_unsigned( 222,8)),
			2470 => std_logic_vector(to_unsigned( 166,8)),
			2471 => std_logic_vector(to_unsigned( 250,8)),
			2472 => std_logic_vector(to_unsigned( 157,8)),
			2473 => std_logic_vector(to_unsigned( 129,8)),
			2474 => std_logic_vector(to_unsigned( 84,8)),
			2475 => std_logic_vector(to_unsigned( 219,8)),
			2476 => std_logic_vector(to_unsigned( 15,8)),
			2477 => std_logic_vector(to_unsigned( 32,8)),
			2478 => std_logic_vector(to_unsigned( 165,8)),
			2479 => std_logic_vector(to_unsigned( 166,8)),
			2480 => std_logic_vector(to_unsigned( 219,8)),
			2481 => std_logic_vector(to_unsigned( 255,8)),
			2482 => std_logic_vector(to_unsigned( 77,8)),
			2483 => std_logic_vector(to_unsigned( 143,8)),
			2484 => std_logic_vector(to_unsigned( 97,8)),
			2485 => std_logic_vector(to_unsigned( 62,8)),
			2486 => std_logic_vector(to_unsigned( 254,8)),
			2487 => std_logic_vector(to_unsigned( 118,8)),
			2488 => std_logic_vector(to_unsigned( 17,8)),
			2489 => std_logic_vector(to_unsigned( 4,8)),
			2490 => std_logic_vector(to_unsigned( 170,8)),
			2491 => std_logic_vector(to_unsigned( 226,8)),
			2492 => std_logic_vector(to_unsigned( 122,8)),
			2493 => std_logic_vector(to_unsigned( 58,8)),
			2494 => std_logic_vector(to_unsigned( 111,8)),
			2495 => std_logic_vector(to_unsigned( 186,8)),
			2496 => std_logic_vector(to_unsigned( 63,8)),
			2497 => std_logic_vector(to_unsigned( 115,8)),
			2498 => std_logic_vector(to_unsigned( 33,8)),
			2499 => std_logic_vector(to_unsigned( 163,8)),
			2500 => std_logic_vector(to_unsigned( 97,8)),
			2501 => std_logic_vector(to_unsigned( 164,8)),
			2502 => std_logic_vector(to_unsigned( 48,8)),
			2503 => std_logic_vector(to_unsigned( 217,8)),
			2504 => std_logic_vector(to_unsigned( 103,8)),
			2505 => std_logic_vector(to_unsigned( 98,8)),
			2506 => std_logic_vector(to_unsigned( 251,8)),
			2507 => std_logic_vector(to_unsigned( 218,8)),
			2508 => std_logic_vector(to_unsigned( 17,8)),
			2509 => std_logic_vector(to_unsigned( 129,8)),
			2510 => std_logic_vector(to_unsigned( 71,8)),
			2511 => std_logic_vector(to_unsigned( 134,8)),
			2512 => std_logic_vector(to_unsigned( 255,8)),
			2513 => std_logic_vector(to_unsigned( 23,8)),
			2514 => std_logic_vector(to_unsigned( 76,8)),
			2515 => std_logic_vector(to_unsigned( 236,8)),
			2516 => std_logic_vector(to_unsigned( 175,8)),
			2517 => std_logic_vector(to_unsigned( 56,8)),
			2518 => std_logic_vector(to_unsigned( 132,8)),
			2519 => std_logic_vector(to_unsigned( 226,8)),
			2520 => std_logic_vector(to_unsigned( 4,8)),
			2521 => std_logic_vector(to_unsigned( 142,8)),
			2522 => std_logic_vector(to_unsigned( 12,8)),
			2523 => std_logic_vector(to_unsigned( 133,8)),
			2524 => std_logic_vector(to_unsigned( 240,8)),
			2525 => std_logic_vector(to_unsigned( 21,8)),
			2526 => std_logic_vector(to_unsigned( 159,8)),
			2527 => std_logic_vector(to_unsigned( 112,8)),
			2528 => std_logic_vector(to_unsigned( 80,8)),
			2529 => std_logic_vector(to_unsigned( 145,8)),
			2530 => std_logic_vector(to_unsigned( 71,8)),
			2531 => std_logic_vector(to_unsigned( 156,8)),
			2532 => std_logic_vector(to_unsigned( 107,8)),
			2533 => std_logic_vector(to_unsigned( 88,8)),
			2534 => std_logic_vector(to_unsigned( 171,8)),
			2535 => std_logic_vector(to_unsigned( 11,8)),
			2536 => std_logic_vector(to_unsigned( 134,8)),
			2537 => std_logic_vector(to_unsigned( 165,8)),
			2538 => std_logic_vector(to_unsigned( 129,8)),
			2539 => std_logic_vector(to_unsigned( 201,8)),
			2540 => std_logic_vector(to_unsigned( 220,8)),
			2541 => std_logic_vector(to_unsigned( 145,8)),
			2542 => std_logic_vector(to_unsigned( 148,8)),
			2543 => std_logic_vector(to_unsigned( 134,8)),
			2544 => std_logic_vector(to_unsigned( 249,8)),
			2545 => std_logic_vector(to_unsigned( 89,8)),
			2546 => std_logic_vector(to_unsigned( 242,8)),
			2547 => std_logic_vector(to_unsigned( 140,8)),
			2548 => std_logic_vector(to_unsigned( 154,8)),
			2549 => std_logic_vector(to_unsigned( 74,8)),
			2550 => std_logic_vector(to_unsigned( 55,8)),
			2551 => std_logic_vector(to_unsigned( 90,8)),
			2552 => std_logic_vector(to_unsigned( 47,8)),
			2553 => std_logic_vector(to_unsigned( 246,8)),
			2554 => std_logic_vector(to_unsigned( 141,8)),
			2555 => std_logic_vector(to_unsigned( 225,8)),
			2556 => std_logic_vector(to_unsigned( 25,8)),
			2557 => std_logic_vector(to_unsigned( 55,8)),
			2558 => std_logic_vector(to_unsigned( 67,8)),
			2559 => std_logic_vector(to_unsigned( 23,8)),
			2560 => std_logic_vector(to_unsigned( 20,8)),
			2561 => std_logic_vector(to_unsigned( 99,8)),
			2562 => std_logic_vector(to_unsigned( 23,8)),
			2563 => std_logic_vector(to_unsigned( 86,8)),
			2564 => std_logic_vector(to_unsigned( 52,8)),
			2565 => std_logic_vector(to_unsigned( 124,8)),
			2566 => std_logic_vector(to_unsigned( 31,8)),
			2567 => std_logic_vector(to_unsigned( 71,8)),
			2568 => std_logic_vector(to_unsigned( 97,8)),
			2569 => std_logic_vector(to_unsigned( 170,8)),
			2570 => std_logic_vector(to_unsigned( 139,8)),
			2571 => std_logic_vector(to_unsigned( 246,8)),
			2572 => std_logic_vector(to_unsigned( 184,8)),
			2573 => std_logic_vector(to_unsigned( 183,8)),
			2574 => std_logic_vector(to_unsigned( 223,8)),
			2575 => std_logic_vector(to_unsigned( 126,8)),
			2576 => std_logic_vector(to_unsigned( 125,8)),
			2577 => std_logic_vector(to_unsigned( 101,8)),
			2578 => std_logic_vector(to_unsigned( 112,8)),
			2579 => std_logic_vector(to_unsigned( 181,8)),
			2580 => std_logic_vector(to_unsigned( 134,8)),
			2581 => std_logic_vector(to_unsigned( 83,8)),
			2582 => std_logic_vector(to_unsigned( 61,8)),
			2583 => std_logic_vector(to_unsigned( 187,8)),
			2584 => std_logic_vector(to_unsigned( 11,8)),
			2585 => std_logic_vector(to_unsigned( 47,8)),
			2586 => std_logic_vector(to_unsigned( 187,8)),
			2587 => std_logic_vector(to_unsigned( 180,8)),
			2588 => std_logic_vector(to_unsigned( 94,8)),
			2589 => std_logic_vector(to_unsigned( 115,8)),
			2590 => std_logic_vector(to_unsigned( 35,8)),
			2591 => std_logic_vector(to_unsigned( 120,8)),
			2592 => std_logic_vector(to_unsigned( 169,8)),
			2593 => std_logic_vector(to_unsigned( 102,8)),
			2594 => std_logic_vector(to_unsigned( 178,8)),
			2595 => std_logic_vector(to_unsigned( 214,8)),
			2596 => std_logic_vector(to_unsigned( 189,8)),
			2597 => std_logic_vector(to_unsigned( 134,8)),
			2598 => std_logic_vector(to_unsigned( 210,8)),
			2599 => std_logic_vector(to_unsigned( 234,8)),
			2600 => std_logic_vector(to_unsigned( 60,8)),
			2601 => std_logic_vector(to_unsigned( 241,8)),
			2602 => std_logic_vector(to_unsigned( 53,8)),
			2603 => std_logic_vector(to_unsigned( 133,8)),
			2604 => std_logic_vector(to_unsigned( 244,8)),
			2605 => std_logic_vector(to_unsigned( 20,8)),
			2606 => std_logic_vector(to_unsigned( 190,8)),
			2607 => std_logic_vector(to_unsigned( 193,8)),
			2608 => std_logic_vector(to_unsigned( 146,8)),
			2609 => std_logic_vector(to_unsigned( 226,8)),
			2610 => std_logic_vector(to_unsigned( 202,8)),
			2611 => std_logic_vector(to_unsigned( 20,8)),
			2612 => std_logic_vector(to_unsigned( 113,8)),
			2613 => std_logic_vector(to_unsigned( 253,8)),
			2614 => std_logic_vector(to_unsigned( 184,8)),
			2615 => std_logic_vector(to_unsigned( 4,8)),
			2616 => std_logic_vector(to_unsigned( 27,8)),
			2617 => std_logic_vector(to_unsigned( 181,8)),
			2618 => std_logic_vector(to_unsigned( 139,8)),
			2619 => std_logic_vector(to_unsigned( 201,8)),
			2620 => std_logic_vector(to_unsigned( 236,8)),
			2621 => std_logic_vector(to_unsigned( 79,8)),
			2622 => std_logic_vector(to_unsigned( 225,8)),
			2623 => std_logic_vector(to_unsigned( 253,8)),
			2624 => std_logic_vector(to_unsigned( 52,8)),
			2625 => std_logic_vector(to_unsigned( 169,8)),
			2626 => std_logic_vector(to_unsigned( 117,8)),
			2627 => std_logic_vector(to_unsigned( 62,8)),
			2628 => std_logic_vector(to_unsigned( 81,8)),
			2629 => std_logic_vector(to_unsigned( 49,8)),
			2630 => std_logic_vector(to_unsigned( 246,8)),
			2631 => std_logic_vector(to_unsigned( 216,8)),
			2632 => std_logic_vector(to_unsigned( 205,8)),
			2633 => std_logic_vector(to_unsigned( 4,8)),
			2634 => std_logic_vector(to_unsigned( 69,8)),
			2635 => std_logic_vector(to_unsigned( 179,8)),
			2636 => std_logic_vector(to_unsigned( 218,8)),
			2637 => std_logic_vector(to_unsigned( 61,8)),
			2638 => std_logic_vector(to_unsigned( 56,8)),
			2639 => std_logic_vector(to_unsigned( 146,8)),
			2640 => std_logic_vector(to_unsigned( 185,8)),
			2641 => std_logic_vector(to_unsigned( 87,8)),
			2642 => std_logic_vector(to_unsigned( 168,8)),
			2643 => std_logic_vector(to_unsigned( 198,8)),
			2644 => std_logic_vector(to_unsigned( 79,8)),
			2645 => std_logic_vector(to_unsigned( 83,8)),
			2646 => std_logic_vector(to_unsigned( 7,8)),
			2647 => std_logic_vector(to_unsigned( 83,8)),
			2648 => std_logic_vector(to_unsigned( 90,8)),
			2649 => std_logic_vector(to_unsigned( 236,8)),
			2650 => std_logic_vector(to_unsigned( 248,8)),
			2651 => std_logic_vector(to_unsigned( 157,8)),
			2652 => std_logic_vector(to_unsigned( 224,8)),
			2653 => std_logic_vector(to_unsigned( 6,8)),
			2654 => std_logic_vector(to_unsigned( 233,8)),
			2655 => std_logic_vector(to_unsigned( 63,8)),
			2656 => std_logic_vector(to_unsigned( 99,8)),
			2657 => std_logic_vector(to_unsigned( 195,8)),
			2658 => std_logic_vector(to_unsigned( 135,8)),
			2659 => std_logic_vector(to_unsigned( 204,8)),
			2660 => std_logic_vector(to_unsigned( 212,8)),
			2661 => std_logic_vector(to_unsigned( 228,8)),
			2662 => std_logic_vector(to_unsigned( 140,8)),
			2663 => std_logic_vector(to_unsigned( 107,8)),
			2664 => std_logic_vector(to_unsigned( 43,8)),
			2665 => std_logic_vector(to_unsigned( 72,8)),
			2666 => std_logic_vector(to_unsigned( 186,8)),
			2667 => std_logic_vector(to_unsigned( 96,8)),
			2668 => std_logic_vector(to_unsigned( 38,8)),
			2669 => std_logic_vector(to_unsigned( 109,8)),
			2670 => std_logic_vector(to_unsigned( 162,8)),
			2671 => std_logic_vector(to_unsigned( 35,8)),
			2672 => std_logic_vector(to_unsigned( 236,8)),
			2673 => std_logic_vector(to_unsigned( 137,8)),
			2674 => std_logic_vector(to_unsigned( 99,8)),
			2675 => std_logic_vector(to_unsigned( 124,8)),
			2676 => std_logic_vector(to_unsigned( 54,8)),
			2677 => std_logic_vector(to_unsigned( 57,8)),
			2678 => std_logic_vector(to_unsigned( 129,8)),
			2679 => std_logic_vector(to_unsigned( 7,8)),
			2680 => std_logic_vector(to_unsigned( 84,8)),
			2681 => std_logic_vector(to_unsigned( 104,8)),
			2682 => std_logic_vector(to_unsigned( 251,8)),
			2683 => std_logic_vector(to_unsigned( 152,8)),
			2684 => std_logic_vector(to_unsigned( 74,8)),
			2685 => std_logic_vector(to_unsigned( 121,8)),
			2686 => std_logic_vector(to_unsigned( 207,8)),
			2687 => std_logic_vector(to_unsigned( 39,8)),
			2688 => std_logic_vector(to_unsigned( 36,8)),
			2689 => std_logic_vector(to_unsigned( 39,8)),
			2690 => std_logic_vector(to_unsigned( 129,8)),
			2691 => std_logic_vector(to_unsigned( 32,8)),
			2692 => std_logic_vector(to_unsigned( 79,8)),
			2693 => std_logic_vector(to_unsigned( 170,8)),
			2694 => std_logic_vector(to_unsigned( 42,8)),
			2695 => std_logic_vector(to_unsigned( 241,8)),
			2696 => std_logic_vector(to_unsigned( 43,8)),
			2697 => std_logic_vector(to_unsigned( 54,8)),
			2698 => std_logic_vector(to_unsigned( 136,8)),
			2699 => std_logic_vector(to_unsigned( 189,8)),
			2700 => std_logic_vector(to_unsigned( 241,8)),
			2701 => std_logic_vector(to_unsigned( 146,8)),
			2702 => std_logic_vector(to_unsigned( 170,8)),
			2703 => std_logic_vector(to_unsigned( 11,8)),
			2704 => std_logic_vector(to_unsigned( 231,8)),
			2705 => std_logic_vector(to_unsigned( 82,8)),
			2706 => std_logic_vector(to_unsigned( 79,8)),
			2707 => std_logic_vector(to_unsigned( 113,8)),
			2708 => std_logic_vector(to_unsigned( 48,8)),
			2709 => std_logic_vector(to_unsigned( 134,8)),
			2710 => std_logic_vector(to_unsigned( 15,8)),
			2711 => std_logic_vector(to_unsigned( 10,8)),
			2712 => std_logic_vector(to_unsigned( 189,8)),
			2713 => std_logic_vector(to_unsigned( 46,8)),
			2714 => std_logic_vector(to_unsigned( 21,8)),
			2715 => std_logic_vector(to_unsigned( 30,8)),
			2716 => std_logic_vector(to_unsigned( 44,8)),
			2717 => std_logic_vector(to_unsigned( 205,8)),
			2718 => std_logic_vector(to_unsigned( 97,8)),
			2719 => std_logic_vector(to_unsigned( 164,8)),
			2720 => std_logic_vector(to_unsigned( 215,8)),
			2721 => std_logic_vector(to_unsigned( 75,8)),
			2722 => std_logic_vector(to_unsigned( 240,8)),
			2723 => std_logic_vector(to_unsigned( 2,8)),
			2724 => std_logic_vector(to_unsigned( 70,8)),
			2725 => std_logic_vector(to_unsigned( 34,8)),
			2726 => std_logic_vector(to_unsigned( 92,8)),
			2727 => std_logic_vector(to_unsigned( 128,8)),
			2728 => std_logic_vector(to_unsigned( 160,8)),
			2729 => std_logic_vector(to_unsigned( 89,8)),
			2730 => std_logic_vector(to_unsigned( 80,8)),
			2731 => std_logic_vector(to_unsigned( 94,8)),
			2732 => std_logic_vector(to_unsigned( 201,8)),
			2733 => std_logic_vector(to_unsigned( 221,8)),
			2734 => std_logic_vector(to_unsigned( 132,8)),
			2735 => std_logic_vector(to_unsigned( 140,8)),
			2736 => std_logic_vector(to_unsigned( 33,8)),
			2737 => std_logic_vector(to_unsigned( 240,8)),
			2738 => std_logic_vector(to_unsigned( 121,8)),
			2739 => std_logic_vector(to_unsigned( 24,8)),
			2740 => std_logic_vector(to_unsigned( 238,8)),
			2741 => std_logic_vector(to_unsigned( 128,8)),
			2742 => std_logic_vector(to_unsigned( 192,8)),
			2743 => std_logic_vector(to_unsigned( 74,8)),
			2744 => std_logic_vector(to_unsigned( 243,8)),
			2745 => std_logic_vector(to_unsigned( 187,8)),
			2746 => std_logic_vector(to_unsigned( 235,8)),
			2747 => std_logic_vector(to_unsigned( 47,8)),
			2748 => std_logic_vector(to_unsigned( 55,8)),
			2749 => std_logic_vector(to_unsigned( 77,8)),
			2750 => std_logic_vector(to_unsigned( 8,8)),
			2751 => std_logic_vector(to_unsigned( 208,8)),
			2752 => std_logic_vector(to_unsigned( 139,8)),
			2753 => std_logic_vector(to_unsigned( 52,8)),
			2754 => std_logic_vector(to_unsigned( 174,8)),
			2755 => std_logic_vector(to_unsigned( 35,8)),
			2756 => std_logic_vector(to_unsigned( 209,8)),
			2757 => std_logic_vector(to_unsigned( 160,8)),
			2758 => std_logic_vector(to_unsigned( 147,8)),
			2759 => std_logic_vector(to_unsigned( 1,8)),
			2760 => std_logic_vector(to_unsigned( 195,8)),
			2761 => std_logic_vector(to_unsigned( 251,8)),
			2762 => std_logic_vector(to_unsigned( 86,8)),
			2763 => std_logic_vector(to_unsigned( 148,8)),
			2764 => std_logic_vector(to_unsigned( 15,8)),
			2765 => std_logic_vector(to_unsigned( 2,8)),
			2766 => std_logic_vector(to_unsigned( 147,8)),
			2767 => std_logic_vector(to_unsigned( 86,8)),
			2768 => std_logic_vector(to_unsigned( 155,8)),
			2769 => std_logic_vector(to_unsigned( 214,8)),
			2770 => std_logic_vector(to_unsigned( 159,8)),
			2771 => std_logic_vector(to_unsigned( 210,8)),
			2772 => std_logic_vector(to_unsigned( 95,8)),
			2773 => std_logic_vector(to_unsigned( 248,8)),
			2774 => std_logic_vector(to_unsigned( 227,8)),
			2775 => std_logic_vector(to_unsigned( 114,8)),
			2776 => std_logic_vector(to_unsigned( 135,8)),
			2777 => std_logic_vector(to_unsigned( 225,8)),
			2778 => std_logic_vector(to_unsigned( 195,8)),
			2779 => std_logic_vector(to_unsigned( 179,8)),
			2780 => std_logic_vector(to_unsigned( 40,8)),
			2781 => std_logic_vector(to_unsigned( 54,8)),
			2782 => std_logic_vector(to_unsigned( 181,8)),
			2783 => std_logic_vector(to_unsigned( 5,8)),
			2784 => std_logic_vector(to_unsigned( 188,8)),
			2785 => std_logic_vector(to_unsigned( 135,8)),
			2786 => std_logic_vector(to_unsigned( 186,8)),
			2787 => std_logic_vector(to_unsigned( 119,8)),
			2788 => std_logic_vector(to_unsigned( 4,8)),
			2789 => std_logic_vector(to_unsigned( 23,8)),
			2790 => std_logic_vector(to_unsigned( 151,8)),
			2791 => std_logic_vector(to_unsigned( 106,8)),
			2792 => std_logic_vector(to_unsigned( 108,8)),
			2793 => std_logic_vector(to_unsigned( 63,8)),
			2794 => std_logic_vector(to_unsigned( 92,8)),
			2795 => std_logic_vector(to_unsigned( 254,8)),
			2796 => std_logic_vector(to_unsigned( 121,8)),
			2797 => std_logic_vector(to_unsigned( 190,8)),
			2798 => std_logic_vector(to_unsigned( 111,8)),
			2799 => std_logic_vector(to_unsigned( 193,8)),
			2800 => std_logic_vector(to_unsigned( 169,8)),
			2801 => std_logic_vector(to_unsigned( 215,8)),
			2802 => std_logic_vector(to_unsigned( 29,8)),
			2803 => std_logic_vector(to_unsigned( 83,8)),
			2804 => std_logic_vector(to_unsigned( 131,8)),
			2805 => std_logic_vector(to_unsigned( 26,8)),
			2806 => std_logic_vector(to_unsigned( 206,8)),
			2807 => std_logic_vector(to_unsigned( 204,8)),
			2808 => std_logic_vector(to_unsigned( 164,8)),
			2809 => std_logic_vector(to_unsigned( 91,8)),
			2810 => std_logic_vector(to_unsigned( 231,8)),
			2811 => std_logic_vector(to_unsigned( 205,8)),
			2812 => std_logic_vector(to_unsigned( 17,8)),
			2813 => std_logic_vector(to_unsigned( 148,8)),
			2814 => std_logic_vector(to_unsigned( 59,8)),
			2815 => std_logic_vector(to_unsigned( 201,8)),
			2816 => std_logic_vector(to_unsigned( 134,8)),
			2817 => std_logic_vector(to_unsigned( 117,8)),
			2818 => std_logic_vector(to_unsigned( 228,8)),
			2819 => std_logic_vector(to_unsigned( 22,8)),
			2820 => std_logic_vector(to_unsigned( 80,8)),
			2821 => std_logic_vector(to_unsigned( 99,8)),
			2822 => std_logic_vector(to_unsigned( 101,8)),
			2823 => std_logic_vector(to_unsigned( 173,8)),
			2824 => std_logic_vector(to_unsigned( 70,8)),
			2825 => std_logic_vector(to_unsigned( 229,8)),
			2826 => std_logic_vector(to_unsigned( 98,8)),
			2827 => std_logic_vector(to_unsigned( 252,8)),
			2828 => std_logic_vector(to_unsigned( 202,8)),
			2829 => std_logic_vector(to_unsigned( 174,8)),
			2830 => std_logic_vector(to_unsigned( 234,8)),
			2831 => std_logic_vector(to_unsigned( 200,8)),
			2832 => std_logic_vector(to_unsigned( 246,8)),
			2833 => std_logic_vector(to_unsigned( 59,8)),
			2834 => std_logic_vector(to_unsigned( 88,8)),
			2835 => std_logic_vector(to_unsigned( 7,8)),
			2836 => std_logic_vector(to_unsigned( 29,8)),
			2837 => std_logic_vector(to_unsigned( 17,8)),
			2838 => std_logic_vector(to_unsigned( 64,8)),
			2839 => std_logic_vector(to_unsigned( 122,8)),
			2840 => std_logic_vector(to_unsigned( 97,8)),
			2841 => std_logic_vector(to_unsigned( 176,8)),
			2842 => std_logic_vector(to_unsigned( 77,8)),
			2843 => std_logic_vector(to_unsigned( 75,8)),
			2844 => std_logic_vector(to_unsigned( 55,8)),
			2845 => std_logic_vector(to_unsigned( 135,8)),
			2846 => std_logic_vector(to_unsigned( 233,8)),
			2847 => std_logic_vector(to_unsigned( 238,8)),
			2848 => std_logic_vector(to_unsigned( 120,8)),
			2849 => std_logic_vector(to_unsigned( 47,8)),
			2850 => std_logic_vector(to_unsigned( 103,8)),
			2851 => std_logic_vector(to_unsigned( 17,8)),
			2852 => std_logic_vector(to_unsigned( 32,8)),
			2853 => std_logic_vector(to_unsigned( 214,8)),
			2854 => std_logic_vector(to_unsigned( 176,8)),
			2855 => std_logic_vector(to_unsigned( 57,8)),
			2856 => std_logic_vector(to_unsigned( 239,8)),
			2857 => std_logic_vector(to_unsigned( 205,8)),
			2858 => std_logic_vector(to_unsigned( 42,8)),
			2859 => std_logic_vector(to_unsigned( 56,8)),
			2860 => std_logic_vector(to_unsigned( 198,8)),
			2861 => std_logic_vector(to_unsigned( 209,8)),
			2862 => std_logic_vector(to_unsigned( 38,8)),
			2863 => std_logic_vector(to_unsigned( 12,8)),
			2864 => std_logic_vector(to_unsigned( 14,8)),
			2865 => std_logic_vector(to_unsigned( 211,8)),
			2866 => std_logic_vector(to_unsigned( 71,8)),
			2867 => std_logic_vector(to_unsigned( 35,8)),
			2868 => std_logic_vector(to_unsigned( 69,8)),
			2869 => std_logic_vector(to_unsigned( 155,8)),
			2870 => std_logic_vector(to_unsigned( 116,8)),
			2871 => std_logic_vector(to_unsigned( 81,8)),
			2872 => std_logic_vector(to_unsigned( 236,8)),
			2873 => std_logic_vector(to_unsigned( 24,8)),
			2874 => std_logic_vector(to_unsigned( 184,8)),
			2875 => std_logic_vector(to_unsigned( 226,8)),
			2876 => std_logic_vector(to_unsigned( 248,8)),
			2877 => std_logic_vector(to_unsigned( 47,8)),
			2878 => std_logic_vector(to_unsigned( 180,8)),
			2879 => std_logic_vector(to_unsigned( 15,8)),
			2880 => std_logic_vector(to_unsigned( 127,8)),
			2881 => std_logic_vector(to_unsigned( 170,8)),
			2882 => std_logic_vector(to_unsigned( 60,8)),
			2883 => std_logic_vector(to_unsigned( 17,8)),
			2884 => std_logic_vector(to_unsigned( 79,8)),
			2885 => std_logic_vector(to_unsigned( 112,8)),
			2886 => std_logic_vector(to_unsigned( 196,8)),
			2887 => std_logic_vector(to_unsigned( 15,8)),
			2888 => std_logic_vector(to_unsigned( 11,8)),
			2889 => std_logic_vector(to_unsigned( 103,8)),
			2890 => std_logic_vector(to_unsigned( 165,8)),
			2891 => std_logic_vector(to_unsigned( 148,8)),
			2892 => std_logic_vector(to_unsigned( 31,8)),
			2893 => std_logic_vector(to_unsigned( 61,8)),
			2894 => std_logic_vector(to_unsigned( 31,8)),
			2895 => std_logic_vector(to_unsigned( 222,8)),
			2896 => std_logic_vector(to_unsigned( 111,8)),
			2897 => std_logic_vector(to_unsigned( 94,8)),
			2898 => std_logic_vector(to_unsigned( 25,8)),
			2899 => std_logic_vector(to_unsigned( 147,8)),
			2900 => std_logic_vector(to_unsigned( 110,8)),
			2901 => std_logic_vector(to_unsigned( 131,8)),
			2902 => std_logic_vector(to_unsigned( 10,8)),
			2903 => std_logic_vector(to_unsigned( 143,8)),
			2904 => std_logic_vector(to_unsigned( 19,8)),
			2905 => std_logic_vector(to_unsigned( 58,8)),
			2906 => std_logic_vector(to_unsigned( 10,8)),
			2907 => std_logic_vector(to_unsigned( 113,8)),
			2908 => std_logic_vector(to_unsigned( 69,8)),
			2909 => std_logic_vector(to_unsigned( 211,8)),
			2910 => std_logic_vector(to_unsigned( 230,8)),
			2911 => std_logic_vector(to_unsigned( 152,8)),
			2912 => std_logic_vector(to_unsigned( 164,8)),
			2913 => std_logic_vector(to_unsigned( 182,8)),
			2914 => std_logic_vector(to_unsigned( 17,8)),
			2915 => std_logic_vector(to_unsigned( 69,8)),
			2916 => std_logic_vector(to_unsigned( 186,8)),
			2917 => std_logic_vector(to_unsigned( 161,8)),
			2918 => std_logic_vector(to_unsigned( 253,8)),
			2919 => std_logic_vector(to_unsigned( 109,8)),
			2920 => std_logic_vector(to_unsigned( 237,8)),
			2921 => std_logic_vector(to_unsigned( 199,8)),
			2922 => std_logic_vector(to_unsigned( 193,8)),
			2923 => std_logic_vector(to_unsigned( 5,8)),
			2924 => std_logic_vector(to_unsigned( 249,8)),
			2925 => std_logic_vector(to_unsigned( 43,8)),
			2926 => std_logic_vector(to_unsigned( 98,8)),
			2927 => std_logic_vector(to_unsigned( 13,8)),
			2928 => std_logic_vector(to_unsigned( 209,8)),
			2929 => std_logic_vector(to_unsigned( 149,8)),
			2930 => std_logic_vector(to_unsigned( 97,8)),
			2931 => std_logic_vector(to_unsigned( 201,8)),
			2932 => std_logic_vector(to_unsigned( 249,8)),
			2933 => std_logic_vector(to_unsigned( 222,8)),
			2934 => std_logic_vector(to_unsigned( 248,8)),
			2935 => std_logic_vector(to_unsigned( 81,8)),
			2936 => std_logic_vector(to_unsigned( 219,8)),
			2937 => std_logic_vector(to_unsigned( 27,8)),
			2938 => std_logic_vector(to_unsigned( 39,8)),
			2939 => std_logic_vector(to_unsigned( 189,8)),
			2940 => std_logic_vector(to_unsigned( 109,8)),
			2941 => std_logic_vector(to_unsigned( 130,8)),
			2942 => std_logic_vector(to_unsigned( 100,8)),
			2943 => std_logic_vector(to_unsigned( 133,8)),
			2944 => std_logic_vector(to_unsigned( 164,8)),
			2945 => std_logic_vector(to_unsigned( 205,8)),
			2946 => std_logic_vector(to_unsigned( 197,8)),
			2947 => std_logic_vector(to_unsigned( 197,8)),
			2948 => std_logic_vector(to_unsigned( 233,8)),
			2949 => std_logic_vector(to_unsigned( 36,8)),
			2950 => std_logic_vector(to_unsigned( 44,8)),
			2951 => std_logic_vector(to_unsigned( 68,8)),
			2952 => std_logic_vector(to_unsigned( 105,8)),
			2953 => std_logic_vector(to_unsigned( 235,8)),
			2954 => std_logic_vector(to_unsigned( 52,8)),
			2955 => std_logic_vector(to_unsigned( 153,8)),
			2956 => std_logic_vector(to_unsigned( 229,8)),
			2957 => std_logic_vector(to_unsigned( 195,8)),
			2958 => std_logic_vector(to_unsigned( 116,8)),
			2959 => std_logic_vector(to_unsigned( 147,8)),
			2960 => std_logic_vector(to_unsigned( 134,8)),
			2961 => std_logic_vector(to_unsigned( 238,8)),
			2962 => std_logic_vector(to_unsigned( 231,8)),
			2963 => std_logic_vector(to_unsigned( 150,8)),
			2964 => std_logic_vector(to_unsigned( 134,8)),
			2965 => std_logic_vector(to_unsigned( 95,8)),
			2966 => std_logic_vector(to_unsigned( 66,8)),
			2967 => std_logic_vector(to_unsigned( 43,8)),
			2968 => std_logic_vector(to_unsigned( 58,8)),
			2969 => std_logic_vector(to_unsigned( 224,8)),
			2970 => std_logic_vector(to_unsigned( 128,8)),
			2971 => std_logic_vector(to_unsigned( 151,8)),
			2972 => std_logic_vector(to_unsigned( 15,8)),
			2973 => std_logic_vector(to_unsigned( 98,8)),
			2974 => std_logic_vector(to_unsigned( 159,8)),
			2975 => std_logic_vector(to_unsigned( 177,8)),
			2976 => std_logic_vector(to_unsigned( 123,8)),
			2977 => std_logic_vector(to_unsigned( 68,8)),
			2978 => std_logic_vector(to_unsigned( 148,8)),
			2979 => std_logic_vector(to_unsigned( 72,8)),
			2980 => std_logic_vector(to_unsigned( 219,8)),
			2981 => std_logic_vector(to_unsigned( 40,8)),
			2982 => std_logic_vector(to_unsigned( 161,8)),
			2983 => std_logic_vector(to_unsigned( 11,8)),
			2984 => std_logic_vector(to_unsigned( 154,8)),
			2985 => std_logic_vector(to_unsigned( 204,8)),
			2986 => std_logic_vector(to_unsigned( 227,8)),
			2987 => std_logic_vector(to_unsigned( 25,8)),
			2988 => std_logic_vector(to_unsigned( 194,8)),
			2989 => std_logic_vector(to_unsigned( 49,8)),
			2990 => std_logic_vector(to_unsigned( 218,8)),
			2991 => std_logic_vector(to_unsigned( 210,8)),
			2992 => std_logic_vector(to_unsigned( 217,8)),
			2993 => std_logic_vector(to_unsigned( 49,8)),
			2994 => std_logic_vector(to_unsigned( 64,8)),
			2995 => std_logic_vector(to_unsigned( 242,8)),
			2996 => std_logic_vector(to_unsigned( 16,8)),
			2997 => std_logic_vector(to_unsigned( 67,8)),
			2998 => std_logic_vector(to_unsigned( 5,8)),
			2999 => std_logic_vector(to_unsigned( 187,8)),
			3000 => std_logic_vector(to_unsigned( 200,8)),
			3001 => std_logic_vector(to_unsigned( 252,8)),
			3002 => std_logic_vector(to_unsigned( 169,8)),
			3003 => std_logic_vector(to_unsigned( 234,8)),
			3004 => std_logic_vector(to_unsigned( 72,8)),
			3005 => std_logic_vector(to_unsigned( 199,8)),
			3006 => std_logic_vector(to_unsigned( 222,8)),
			3007 => std_logic_vector(to_unsigned( 208,8)),
			3008 => std_logic_vector(to_unsigned( 70,8)),
			3009 => std_logic_vector(to_unsigned( 230,8)),
			3010 => std_logic_vector(to_unsigned( 106,8)),
			3011 => std_logic_vector(to_unsigned( 19,8)),
			3012 => std_logic_vector(to_unsigned( 91,8)),
			3013 => std_logic_vector(to_unsigned( 201,8)),
			3014 => std_logic_vector(to_unsigned( 77,8)),
			3015 => std_logic_vector(to_unsigned( 226,8)),
			3016 => std_logic_vector(to_unsigned( 53,8)),
			3017 => std_logic_vector(to_unsigned( 55,8)),
			3018 => std_logic_vector(to_unsigned( 102,8)),
			3019 => std_logic_vector(to_unsigned( 121,8)),
			3020 => std_logic_vector(to_unsigned( 222,8)),
			3021 => std_logic_vector(to_unsigned( 179,8)),
			3022 => std_logic_vector(to_unsigned( 146,8)),
			3023 => std_logic_vector(to_unsigned( 113,8)),
			3024 => std_logic_vector(to_unsigned( 13,8)),
			3025 => std_logic_vector(to_unsigned( 124,8)),
			3026 => std_logic_vector(to_unsigned( 31,8)),
			3027 => std_logic_vector(to_unsigned( 187,8)),
			3028 => std_logic_vector(to_unsigned( 148,8)),
			3029 => std_logic_vector(to_unsigned( 94,8)),
			3030 => std_logic_vector(to_unsigned( 138,8)),
			3031 => std_logic_vector(to_unsigned( 194,8)),
			3032 => std_logic_vector(to_unsigned( 109,8)),
			3033 => std_logic_vector(to_unsigned( 154,8)),
			3034 => std_logic_vector(to_unsigned( 151,8)),
			3035 => std_logic_vector(to_unsigned( 207,8)),
			3036 => std_logic_vector(to_unsigned( 74,8)),
			3037 => std_logic_vector(to_unsigned( 170,8)),
			3038 => std_logic_vector(to_unsigned( 22,8)),
			3039 => std_logic_vector(to_unsigned( 90,8)),
			3040 => std_logic_vector(to_unsigned( 121,8)),
			3041 => std_logic_vector(to_unsigned( 200,8)),
			3042 => std_logic_vector(to_unsigned( 54,8)),
			3043 => std_logic_vector(to_unsigned( 123,8)),
			3044 => std_logic_vector(to_unsigned( 3,8)),
			3045 => std_logic_vector(to_unsigned( 108,8)),
			3046 => std_logic_vector(to_unsigned( 86,8)),
			3047 => std_logic_vector(to_unsigned( 226,8)),
			3048 => std_logic_vector(to_unsigned( 78,8)),
			3049 => std_logic_vector(to_unsigned( 145,8)),
			3050 => std_logic_vector(to_unsigned( 51,8)),
			3051 => std_logic_vector(to_unsigned( 103,8)),
			3052 => std_logic_vector(to_unsigned( 240,8)),
			3053 => std_logic_vector(to_unsigned( 144,8)),
			3054 => std_logic_vector(to_unsigned( 193,8)),
			3055 => std_logic_vector(to_unsigned( 203,8)),
			3056 => std_logic_vector(to_unsigned( 161,8)),
			3057 => std_logic_vector(to_unsigned( 133,8)),
			3058 => std_logic_vector(to_unsigned( 101,8)),
			3059 => std_logic_vector(to_unsigned( 158,8)),
			3060 => std_logic_vector(to_unsigned( 116,8)),
			3061 => std_logic_vector(to_unsigned( 219,8)),
			3062 => std_logic_vector(to_unsigned( 137,8)),
			3063 => std_logic_vector(to_unsigned( 15,8)),
			3064 => std_logic_vector(to_unsigned( 222,8)),
			3065 => std_logic_vector(to_unsigned( 243,8)),
			3066 => std_logic_vector(to_unsigned( 134,8)),
			3067 => std_logic_vector(to_unsigned( 104,8)),
			3068 => std_logic_vector(to_unsigned( 215,8)),
			3069 => std_logic_vector(to_unsigned( 144,8)),
			3070 => std_logic_vector(to_unsigned( 133,8)),
			3071 => std_logic_vector(to_unsigned( 127,8)),
			3072 => std_logic_vector(to_unsigned( 119,8)),
			3073 => std_logic_vector(to_unsigned( 147,8)),
			3074 => std_logic_vector(to_unsigned( 226,8)),
			3075 => std_logic_vector(to_unsigned( 168,8)),
			3076 => std_logic_vector(to_unsigned( 243,8)),
			3077 => std_logic_vector(to_unsigned( 253,8)),
			3078 => std_logic_vector(to_unsigned( 106,8)),
			3079 => std_logic_vector(to_unsigned( 36,8)),
			3080 => std_logic_vector(to_unsigned( 135,8)),
			3081 => std_logic_vector(to_unsigned( 244,8)),
			3082 => std_logic_vector(to_unsigned( 222,8)),
			3083 => std_logic_vector(to_unsigned( 31,8)),
			3084 => std_logic_vector(to_unsigned( 222,8)),
			3085 => std_logic_vector(to_unsigned( 199,8)),
			3086 => std_logic_vector(to_unsigned( 92,8)),
			3087 => std_logic_vector(to_unsigned( 199,8)),
			3088 => std_logic_vector(to_unsigned( 25,8)),
			3089 => std_logic_vector(to_unsigned( 179,8)),
			3090 => std_logic_vector(to_unsigned( 102,8)),
			3091 => std_logic_vector(to_unsigned( 227,8)),
			3092 => std_logic_vector(to_unsigned( 44,8)),
			3093 => std_logic_vector(to_unsigned( 5,8)),
			3094 => std_logic_vector(to_unsigned( 99,8)),
			3095 => std_logic_vector(to_unsigned( 250,8)),
			3096 => std_logic_vector(to_unsigned( 199,8)),
			3097 => std_logic_vector(to_unsigned( 1,8)),
			3098 => std_logic_vector(to_unsigned( 124,8)),
			3099 => std_logic_vector(to_unsigned( 190,8)),
			3100 => std_logic_vector(to_unsigned( 61,8)),
			3101 => std_logic_vector(to_unsigned( 210,8)),
			3102 => std_logic_vector(to_unsigned( 185,8)),
			3103 => std_logic_vector(to_unsigned( 253,8)),
			3104 => std_logic_vector(to_unsigned( 164,8)),
			3105 => std_logic_vector(to_unsigned( 141,8)),
			3106 => std_logic_vector(to_unsigned( 246,8)),
			3107 => std_logic_vector(to_unsigned( 182,8)),
			3108 => std_logic_vector(to_unsigned( 184,8)),
			3109 => std_logic_vector(to_unsigned( 216,8)),
			3110 => std_logic_vector(to_unsigned( 188,8)),
			3111 => std_logic_vector(to_unsigned( 62,8)),
			3112 => std_logic_vector(to_unsigned( 122,8)),
			3113 => std_logic_vector(to_unsigned( 66,8)),
			3114 => std_logic_vector(to_unsigned( 28,8)),
			3115 => std_logic_vector(to_unsigned( 158,8)),
			3116 => std_logic_vector(to_unsigned( 66,8)),
			3117 => std_logic_vector(to_unsigned( 65,8)),
			3118 => std_logic_vector(to_unsigned( 93,8)),
			3119 => std_logic_vector(to_unsigned( 239,8)),
			3120 => std_logic_vector(to_unsigned( 146,8)),
			3121 => std_logic_vector(to_unsigned( 25,8)),
			3122 => std_logic_vector(to_unsigned( 9,8)),
			3123 => std_logic_vector(to_unsigned( 54,8)),
			3124 => std_logic_vector(to_unsigned( 136,8)),
			3125 => std_logic_vector(to_unsigned( 119,8)),
			3126 => std_logic_vector(to_unsigned( 129,8)),
			3127 => std_logic_vector(to_unsigned( 92,8)),
			3128 => std_logic_vector(to_unsigned( 116,8)),
			3129 => std_logic_vector(to_unsigned( 19,8)),
			3130 => std_logic_vector(to_unsigned( 151,8)),
			3131 => std_logic_vector(to_unsigned( 139,8)),
			3132 => std_logic_vector(to_unsigned( 8,8)),
			3133 => std_logic_vector(to_unsigned( 164,8)),
			3134 => std_logic_vector(to_unsigned( 72,8)),
			3135 => std_logic_vector(to_unsigned( 121,8)),
			3136 => std_logic_vector(to_unsigned( 1,8)),
			3137 => std_logic_vector(to_unsigned( 41,8)),
			3138 => std_logic_vector(to_unsigned( 14,8)),
			3139 => std_logic_vector(to_unsigned( 117,8)),
			3140 => std_logic_vector(to_unsigned( 209,8)),
			3141 => std_logic_vector(to_unsigned( 57,8)),
			3142 => std_logic_vector(to_unsigned( 50,8)),
			3143 => std_logic_vector(to_unsigned( 134,8)),
			3144 => std_logic_vector(to_unsigned( 17,8)),
			3145 => std_logic_vector(to_unsigned( 215,8)),
			3146 => std_logic_vector(to_unsigned( 181,8)),
			3147 => std_logic_vector(to_unsigned( 247,8)),
			3148 => std_logic_vector(to_unsigned( 67,8)),
			3149 => std_logic_vector(to_unsigned( 254,8)),
			3150 => std_logic_vector(to_unsigned( 71,8)),
			3151 => std_logic_vector(to_unsigned( 66,8)),
			3152 => std_logic_vector(to_unsigned( 149,8)),
			3153 => std_logic_vector(to_unsigned( 20,8)),
			3154 => std_logic_vector(to_unsigned( 232,8)),
			3155 => std_logic_vector(to_unsigned( 99,8)),
			3156 => std_logic_vector(to_unsigned( 251,8)),
			3157 => std_logic_vector(to_unsigned( 44,8)),
			3158 => std_logic_vector(to_unsigned( 156,8)),
			3159 => std_logic_vector(to_unsigned( 192,8)),
			3160 => std_logic_vector(to_unsigned( 185,8)),
			3161 => std_logic_vector(to_unsigned( 143,8)),
			3162 => std_logic_vector(to_unsigned( 16,8)),
			3163 => std_logic_vector(to_unsigned( 162,8)),
			3164 => std_logic_vector(to_unsigned( 11,8)),
			3165 => std_logic_vector(to_unsigned( 124,8)),
			3166 => std_logic_vector(to_unsigned( 202,8)),
			3167 => std_logic_vector(to_unsigned( 246,8)),
			3168 => std_logic_vector(to_unsigned( 88,8)),
			3169 => std_logic_vector(to_unsigned( 147,8)),
			3170 => std_logic_vector(to_unsigned( 37,8)),
			3171 => std_logic_vector(to_unsigned( 88,8)),
			3172 => std_logic_vector(to_unsigned( 1,8)),
			3173 => std_logic_vector(to_unsigned( 52,8)),
			3174 => std_logic_vector(to_unsigned( 241,8)),
			3175 => std_logic_vector(to_unsigned( 59,8)),
			3176 => std_logic_vector(to_unsigned( 215,8)),
			3177 => std_logic_vector(to_unsigned( 16,8)),
			3178 => std_logic_vector(to_unsigned( 99,8)),
			3179 => std_logic_vector(to_unsigned( 89,8)),
			3180 => std_logic_vector(to_unsigned( 72,8)),
			3181 => std_logic_vector(to_unsigned( 147,8)),
			3182 => std_logic_vector(to_unsigned( 17,8)),
			3183 => std_logic_vector(to_unsigned( 149,8)),
			3184 => std_logic_vector(to_unsigned( 228,8)),
			3185 => std_logic_vector(to_unsigned( 178,8)),
			3186 => std_logic_vector(to_unsigned( 119,8)),
			3187 => std_logic_vector(to_unsigned( 203,8)),
			3188 => std_logic_vector(to_unsigned( 77,8)),
			3189 => std_logic_vector(to_unsigned( 141,8)),
			3190 => std_logic_vector(to_unsigned( 168,8)),
			3191 => std_logic_vector(to_unsigned( 184,8)),
			3192 => std_logic_vector(to_unsigned( 47,8)),
			3193 => std_logic_vector(to_unsigned( 142,8)),
			3194 => std_logic_vector(to_unsigned( 195,8)),
			3195 => std_logic_vector(to_unsigned( 28,8)),
			3196 => std_logic_vector(to_unsigned( 45,8)),
			3197 => std_logic_vector(to_unsigned( 177,8)),
			3198 => std_logic_vector(to_unsigned( 2,8)),
			3199 => std_logic_vector(to_unsigned( 15,8)),
			3200 => std_logic_vector(to_unsigned( 122,8)),
			3201 => std_logic_vector(to_unsigned( 45,8)),
			3202 => std_logic_vector(to_unsigned( 199,8)),
			3203 => std_logic_vector(to_unsigned( 1,8)),
			3204 => std_logic_vector(to_unsigned( 240,8)),
			3205 => std_logic_vector(to_unsigned( 192,8)),
			3206 => std_logic_vector(to_unsigned( 105,8)),
			3207 => std_logic_vector(to_unsigned( 246,8)),
			3208 => std_logic_vector(to_unsigned( 197,8)),
			3209 => std_logic_vector(to_unsigned( 38,8)),
			3210 => std_logic_vector(to_unsigned( 160,8)),
			3211 => std_logic_vector(to_unsigned( 130,8)),
			3212 => std_logic_vector(to_unsigned( 42,8)),
			3213 => std_logic_vector(to_unsigned( 206,8)),
			3214 => std_logic_vector(to_unsigned( 192,8)),
			3215 => std_logic_vector(to_unsigned( 225,8)),
			3216 => std_logic_vector(to_unsigned( 232,8)),
			3217 => std_logic_vector(to_unsigned( 117,8)),
			3218 => std_logic_vector(to_unsigned( 215,8)),
			3219 => std_logic_vector(to_unsigned( 61,8)),
			3220 => std_logic_vector(to_unsigned( 255,8)),
			3221 => std_logic_vector(to_unsigned( 44,8)),
			3222 => std_logic_vector(to_unsigned( 107,8)),
			3223 => std_logic_vector(to_unsigned( 61,8)),
			3224 => std_logic_vector(to_unsigned( 16,8)),
			3225 => std_logic_vector(to_unsigned( 247,8)),
			3226 => std_logic_vector(to_unsigned( 227,8)),
			3227 => std_logic_vector(to_unsigned( 120,8)),
			3228 => std_logic_vector(to_unsigned( 227,8)),
			3229 => std_logic_vector(to_unsigned( 142,8)),
			3230 => std_logic_vector(to_unsigned( 133,8)),
			3231 => std_logic_vector(to_unsigned( 168,8)),
			3232 => std_logic_vector(to_unsigned( 110,8)),
			3233 => std_logic_vector(to_unsigned( 197,8)),
			3234 => std_logic_vector(to_unsigned( 39,8)),
			3235 => std_logic_vector(to_unsigned( 18,8)),
			3236 => std_logic_vector(to_unsigned( 174,8)),
			3237 => std_logic_vector(to_unsigned( 168,8)),
			3238 => std_logic_vector(to_unsigned( 25,8)),
			3239 => std_logic_vector(to_unsigned( 94,8)),
			3240 => std_logic_vector(to_unsigned( 107,8)),
			3241 => std_logic_vector(to_unsigned( 201,8)),
			3242 => std_logic_vector(to_unsigned( 232,8)),
			3243 => std_logic_vector(to_unsigned( 117,8)),
			3244 => std_logic_vector(to_unsigned( 13,8)),
			3245 => std_logic_vector(to_unsigned( 194,8)),
			3246 => std_logic_vector(to_unsigned( 166,8)),
			3247 => std_logic_vector(to_unsigned( 31,8)),
			3248 => std_logic_vector(to_unsigned( 110,8)),
			3249 => std_logic_vector(to_unsigned( 196,8)),
			3250 => std_logic_vector(to_unsigned( 225,8)),
			3251 => std_logic_vector(to_unsigned( 143,8)),
			3252 => std_logic_vector(to_unsigned( 234,8)),
			3253 => std_logic_vector(to_unsigned( 149,8)),
			3254 => std_logic_vector(to_unsigned( 138,8)),
			3255 => std_logic_vector(to_unsigned( 227,8)),
			3256 => std_logic_vector(to_unsigned( 77,8)),
			3257 => std_logic_vector(to_unsigned( 192,8)),
			3258 => std_logic_vector(to_unsigned( 172,8)),
			3259 => std_logic_vector(to_unsigned( 212,8)),
			3260 => std_logic_vector(to_unsigned( 30,8)),
			3261 => std_logic_vector(to_unsigned( 69,8)),
			3262 => std_logic_vector(to_unsigned( 99,8)),
			3263 => std_logic_vector(to_unsigned( 178,8)),
			3264 => std_logic_vector(to_unsigned( 169,8)),
			3265 => std_logic_vector(to_unsigned( 26,8)),
			3266 => std_logic_vector(to_unsigned( 192,8)),
			3267 => std_logic_vector(to_unsigned( 174,8)),
			3268 => std_logic_vector(to_unsigned( 104,8)),
			3269 => std_logic_vector(to_unsigned( 232,8)),
			3270 => std_logic_vector(to_unsigned( 111,8)),
			3271 => std_logic_vector(to_unsigned( 127,8)),
			3272 => std_logic_vector(to_unsigned( 71,8)),
			3273 => std_logic_vector(to_unsigned( 73,8)),
			3274 => std_logic_vector(to_unsigned( 233,8)),
			3275 => std_logic_vector(to_unsigned( 6,8)),
			3276 => std_logic_vector(to_unsigned( 143,8)),
			3277 => std_logic_vector(to_unsigned( 127,8)),
			3278 => std_logic_vector(to_unsigned( 121,8)),
			3279 => std_logic_vector(to_unsigned( 184,8)),
			3280 => std_logic_vector(to_unsigned( 237,8)),
			3281 => std_logic_vector(to_unsigned( 168,8)),
			3282 => std_logic_vector(to_unsigned( 163,8)),
			3283 => std_logic_vector(to_unsigned( 38,8)),
			3284 => std_logic_vector(to_unsigned( 143,8)),
			3285 => std_logic_vector(to_unsigned( 209,8)),
			3286 => std_logic_vector(to_unsigned( 32,8)),
			3287 => std_logic_vector(to_unsigned( 251,8)),
			3288 => std_logic_vector(to_unsigned( 164,8)),
			3289 => std_logic_vector(to_unsigned( 157,8)),
			3290 => std_logic_vector(to_unsigned( 219,8)),
			3291 => std_logic_vector(to_unsigned( 136,8)),
			3292 => std_logic_vector(to_unsigned( 255,8)),
			3293 => std_logic_vector(to_unsigned( 244,8)),
			3294 => std_logic_vector(to_unsigned( 84,8)),
			3295 => std_logic_vector(to_unsigned( 147,8)),
			3296 => std_logic_vector(to_unsigned( 230,8)),
			3297 => std_logic_vector(to_unsigned( 9,8)),
			3298 => std_logic_vector(to_unsigned( 177,8)),
			3299 => std_logic_vector(to_unsigned( 81,8)),
			3300 => std_logic_vector(to_unsigned( 35,8)),
			3301 => std_logic_vector(to_unsigned( 119,8)),
			3302 => std_logic_vector(to_unsigned( 97,8)),
			3303 => std_logic_vector(to_unsigned( 179,8)),
			3304 => std_logic_vector(to_unsigned( 177,8)),
			3305 => std_logic_vector(to_unsigned( 23,8)),
			3306 => std_logic_vector(to_unsigned( 123,8)),
			3307 => std_logic_vector(to_unsigned( 219,8)),
			3308 => std_logic_vector(to_unsigned( 108,8)),
			3309 => std_logic_vector(to_unsigned( 132,8)),
			3310 => std_logic_vector(to_unsigned( 174,8)),
			3311 => std_logic_vector(to_unsigned( 27,8)),
			3312 => std_logic_vector(to_unsigned( 3,8)),
			3313 => std_logic_vector(to_unsigned( 87,8)),
			3314 => std_logic_vector(to_unsigned( 170,8)),
			3315 => std_logic_vector(to_unsigned( 103,8)),
			3316 => std_logic_vector(to_unsigned( 12,8)),
			3317 => std_logic_vector(to_unsigned( 144,8)),
			3318 => std_logic_vector(to_unsigned( 170,8)),
			3319 => std_logic_vector(to_unsigned( 87,8)),
			3320 => std_logic_vector(to_unsigned( 237,8)),
			3321 => std_logic_vector(to_unsigned( 74,8)),
			3322 => std_logic_vector(to_unsigned( 187,8)),
			3323 => std_logic_vector(to_unsigned( 61,8)),
			3324 => std_logic_vector(to_unsigned( 33,8)),
			3325 => std_logic_vector(to_unsigned( 20,8)),
			3326 => std_logic_vector(to_unsigned( 170,8)),
			3327 => std_logic_vector(to_unsigned( 73,8)),
			3328 => std_logic_vector(to_unsigned( 28,8)),
			3329 => std_logic_vector(to_unsigned( 91,8)),
			3330 => std_logic_vector(to_unsigned( 169,8)),
			3331 => std_logic_vector(to_unsigned( 31,8)),
			3332 => std_logic_vector(to_unsigned( 139,8)),
			3333 => std_logic_vector(to_unsigned( 237,8)),
			3334 => std_logic_vector(to_unsigned( 10,8)),
			3335 => std_logic_vector(to_unsigned( 28,8)),
			3336 => std_logic_vector(to_unsigned( 20,8)),
			3337 => std_logic_vector(to_unsigned( 199,8)),
			3338 => std_logic_vector(to_unsigned( 159,8)),
			3339 => std_logic_vector(to_unsigned( 192,8)),
			3340 => std_logic_vector(to_unsigned( 133,8)),
			3341 => std_logic_vector(to_unsigned( 206,8)),
			3342 => std_logic_vector(to_unsigned( 255,8)),
			3343 => std_logic_vector(to_unsigned( 129,8)),
			3344 => std_logic_vector(to_unsigned( 90,8)),
			3345 => std_logic_vector(to_unsigned( 14,8)),
			3346 => std_logic_vector(to_unsigned( 107,8)),
			3347 => std_logic_vector(to_unsigned( 186,8)),
			3348 => std_logic_vector(to_unsigned( 20,8)),
			3349 => std_logic_vector(to_unsigned( 182,8)),
			3350 => std_logic_vector(to_unsigned( 20,8)),
			3351 => std_logic_vector(to_unsigned( 225,8)),
			3352 => std_logic_vector(to_unsigned( 137,8)),
			3353 => std_logic_vector(to_unsigned( 87,8)),
			3354 => std_logic_vector(to_unsigned( 33,8)),
			3355 => std_logic_vector(to_unsigned( 120,8)),
			3356 => std_logic_vector(to_unsigned( 209,8)),
			3357 => std_logic_vector(to_unsigned( 149,8)),
			3358 => std_logic_vector(to_unsigned( 200,8)),
			3359 => std_logic_vector(to_unsigned( 233,8)),
			3360 => std_logic_vector(to_unsigned( 74,8)),
			3361 => std_logic_vector(to_unsigned( 176,8)),
			3362 => std_logic_vector(to_unsigned( 192,8)),
			3363 => std_logic_vector(to_unsigned( 238,8)),
			3364 => std_logic_vector(to_unsigned( 66,8)),
			3365 => std_logic_vector(to_unsigned( 216,8)),
			3366 => std_logic_vector(to_unsigned( 33,8)),
			3367 => std_logic_vector(to_unsigned( 94,8)),
			3368 => std_logic_vector(to_unsigned( 16,8)),
			3369 => std_logic_vector(to_unsigned( 108,8)),
			3370 => std_logic_vector(to_unsigned( 234,8)),
			3371 => std_logic_vector(to_unsigned( 237,8)),
			3372 => std_logic_vector(to_unsigned( 164,8)),
			3373 => std_logic_vector(to_unsigned( 112,8)),
			3374 => std_logic_vector(to_unsigned( 210,8)),
			3375 => std_logic_vector(to_unsigned( 25,8)),
			3376 => std_logic_vector(to_unsigned( 231,8)),
			3377 => std_logic_vector(to_unsigned( 94,8)),
			3378 => std_logic_vector(to_unsigned( 5,8)),
			3379 => std_logic_vector(to_unsigned( 210,8)),
			3380 => std_logic_vector(to_unsigned( 153,8)),
			3381 => std_logic_vector(to_unsigned( 219,8)),
			3382 => std_logic_vector(to_unsigned( 104,8)),
			3383 => std_logic_vector(to_unsigned( 144,8)),
			3384 => std_logic_vector(to_unsigned( 119,8)),
			3385 => std_logic_vector(to_unsigned( 242,8)),
			3386 => std_logic_vector(to_unsigned( 32,8)),
			3387 => std_logic_vector(to_unsigned( 91,8)),
			3388 => std_logic_vector(to_unsigned( 149,8)),
			3389 => std_logic_vector(to_unsigned( 165,8)),
			3390 => std_logic_vector(to_unsigned( 70,8)),
			3391 => std_logic_vector(to_unsigned( 30,8)),
			3392 => std_logic_vector(to_unsigned( 212,8)),
			3393 => std_logic_vector(to_unsigned( 220,8)),
			3394 => std_logic_vector(to_unsigned( 75,8)),
			3395 => std_logic_vector(to_unsigned( 83,8)),
			3396 => std_logic_vector(to_unsigned( 245,8)),
			3397 => std_logic_vector(to_unsigned( 250,8)),
			3398 => std_logic_vector(to_unsigned( 243,8)),
			3399 => std_logic_vector(to_unsigned( 127,8)),
			3400 => std_logic_vector(to_unsigned( 130,8)),
			3401 => std_logic_vector(to_unsigned( 238,8)),
			3402 => std_logic_vector(to_unsigned( 76,8)),
			3403 => std_logic_vector(to_unsigned( 83,8)),
			3404 => std_logic_vector(to_unsigned( 44,8)),
			3405 => std_logic_vector(to_unsigned( 243,8)),
			3406 => std_logic_vector(to_unsigned( 250,8)),
			3407 => std_logic_vector(to_unsigned( 29,8)),
			3408 => std_logic_vector(to_unsigned( 185,8)),
			3409 => std_logic_vector(to_unsigned( 92,8)),
			3410 => std_logic_vector(to_unsigned( 18,8)),
			3411 => std_logic_vector(to_unsigned( 1,8)),
			3412 => std_logic_vector(to_unsigned( 199,8)),
			3413 => std_logic_vector(to_unsigned( 100,8)),
			3414 => std_logic_vector(to_unsigned( 45,8)),
			3415 => std_logic_vector(to_unsigned( 191,8)),
			3416 => std_logic_vector(to_unsigned( 133,8)),
			3417 => std_logic_vector(to_unsigned( 10,8)),
			3418 => std_logic_vector(to_unsigned( 147,8)),
			3419 => std_logic_vector(to_unsigned( 143,8)),
			3420 => std_logic_vector(to_unsigned( 104,8)),
			3421 => std_logic_vector(to_unsigned( 241,8)),
			3422 => std_logic_vector(to_unsigned( 158,8)),
			3423 => std_logic_vector(to_unsigned( 215,8)),
			3424 => std_logic_vector(to_unsigned( 26,8)),
			3425 => std_logic_vector(to_unsigned( 66,8)),
			3426 => std_logic_vector(to_unsigned( 223,8)),
			3427 => std_logic_vector(to_unsigned( 13,8)),
			3428 => std_logic_vector(to_unsigned( 225,8)),
			3429 => std_logic_vector(to_unsigned( 187,8)),
			3430 => std_logic_vector(to_unsigned( 167,8)),
			3431 => std_logic_vector(to_unsigned( 202,8)),
			3432 => std_logic_vector(to_unsigned( 41,8)),
			3433 => std_logic_vector(to_unsigned( 91,8)),
			3434 => std_logic_vector(to_unsigned( 198,8)),
			3435 => std_logic_vector(to_unsigned( 83,8)),
			3436 => std_logic_vector(to_unsigned( 228,8)),
			3437 => std_logic_vector(to_unsigned( 22,8)),
			3438 => std_logic_vector(to_unsigned( 159,8)),
			3439 => std_logic_vector(to_unsigned( 12,8)),
			3440 => std_logic_vector(to_unsigned( 34,8)),
			3441 => std_logic_vector(to_unsigned( 226,8)),
			3442 => std_logic_vector(to_unsigned( 148,8)),
			3443 => std_logic_vector(to_unsigned( 55,8)),
			3444 => std_logic_vector(to_unsigned( 177,8)),
			3445 => std_logic_vector(to_unsigned( 34,8)),
			3446 => std_logic_vector(to_unsigned( 227,8)),
			3447 => std_logic_vector(to_unsigned( 62,8)),
			3448 => std_logic_vector(to_unsigned( 217,8)),
			3449 => std_logic_vector(to_unsigned( 90,8)),
			3450 => std_logic_vector(to_unsigned( 209,8)),
			3451 => std_logic_vector(to_unsigned( 175,8)),
			3452 => std_logic_vector(to_unsigned( 184,8)),
			3453 => std_logic_vector(to_unsigned( 168,8)),
			3454 => std_logic_vector(to_unsigned( 0,8)),
			3455 => std_logic_vector(to_unsigned( 28,8)),
			3456 => std_logic_vector(to_unsigned( 125,8)),
			3457 => std_logic_vector(to_unsigned( 151,8)),
			3458 => std_logic_vector(to_unsigned( 124,8)),
			3459 => std_logic_vector(to_unsigned( 44,8)),
			3460 => std_logic_vector(to_unsigned( 82,8)),
			3461 => std_logic_vector(to_unsigned( 64,8)),
			3462 => std_logic_vector(to_unsigned( 216,8)),
			3463 => std_logic_vector(to_unsigned( 23,8)),
			3464 => std_logic_vector(to_unsigned( 29,8)),
			3465 => std_logic_vector(to_unsigned( 245,8)),
			3466 => std_logic_vector(to_unsigned( 169,8)),
			3467 => std_logic_vector(to_unsigned( 57,8)),
			3468 => std_logic_vector(to_unsigned( 1,8)),
			3469 => std_logic_vector(to_unsigned( 86,8)),
			3470 => std_logic_vector(to_unsigned( 3,8)),
			3471 => std_logic_vector(to_unsigned( 240,8)),
			3472 => std_logic_vector(to_unsigned( 75,8)),
			3473 => std_logic_vector(to_unsigned( 125,8)),
			3474 => std_logic_vector(to_unsigned( 200,8)),
			3475 => std_logic_vector(to_unsigned( 186,8)),
			3476 => std_logic_vector(to_unsigned( 224,8)),
			3477 => std_logic_vector(to_unsigned( 87,8)),
			3478 => std_logic_vector(to_unsigned( 188,8)),
			3479 => std_logic_vector(to_unsigned( 28,8)),
			3480 => std_logic_vector(to_unsigned( 117,8)),
			3481 => std_logic_vector(to_unsigned( 1,8)),
			3482 => std_logic_vector(to_unsigned( 202,8)),
			3483 => std_logic_vector(to_unsigned( 177,8)),
			3484 => std_logic_vector(to_unsigned( 142,8)),
			3485 => std_logic_vector(to_unsigned( 119,8)),
			3486 => std_logic_vector(to_unsigned( 180,8)),
			3487 => std_logic_vector(to_unsigned( 211,8)),
			3488 => std_logic_vector(to_unsigned( 207,8)),
			3489 => std_logic_vector(to_unsigned( 121,8)),
			3490 => std_logic_vector(to_unsigned( 216,8)),
			3491 => std_logic_vector(to_unsigned( 23,8)),
			3492 => std_logic_vector(to_unsigned( 198,8)),
			3493 => std_logic_vector(to_unsigned( 72,8)),
			3494 => std_logic_vector(to_unsigned( 169,8)),
			3495 => std_logic_vector(to_unsigned( 30,8)),
			3496 => std_logic_vector(to_unsigned( 49,8)),
			3497 => std_logic_vector(to_unsigned( 93,8)),
			3498 => std_logic_vector(to_unsigned( 196,8)),
			3499 => std_logic_vector(to_unsigned( 208,8)),
			3500 => std_logic_vector(to_unsigned( 212,8)),
			3501 => std_logic_vector(to_unsigned( 66,8)),
			3502 => std_logic_vector(to_unsigned( 37,8)),
			3503 => std_logic_vector(to_unsigned( 85,8)),
			3504 => std_logic_vector(to_unsigned( 100,8)),
			3505 => std_logic_vector(to_unsigned( 2,8)),
			3506 => std_logic_vector(to_unsigned( 223,8)),
			3507 => std_logic_vector(to_unsigned( 70,8)),
			3508 => std_logic_vector(to_unsigned( 24,8)),
			3509 => std_logic_vector(to_unsigned( 232,8)),
			3510 => std_logic_vector(to_unsigned( 1,8)),
			3511 => std_logic_vector(to_unsigned( 251,8)),
			3512 => std_logic_vector(to_unsigned( 8,8)),
			3513 => std_logic_vector(to_unsigned( 208,8)),
			3514 => std_logic_vector(to_unsigned( 28,8)),
			3515 => std_logic_vector(to_unsigned( 128,8)),
			3516 => std_logic_vector(to_unsigned( 8,8)),
			3517 => std_logic_vector(to_unsigned( 204,8)),
			3518 => std_logic_vector(to_unsigned( 245,8)),
			3519 => std_logic_vector(to_unsigned( 177,8)),
			3520 => std_logic_vector(to_unsigned( 218,8)),
			3521 => std_logic_vector(to_unsigned( 60,8)),
			3522 => std_logic_vector(to_unsigned( 55,8)),
			3523 => std_logic_vector(to_unsigned( 142,8)),
			3524 => std_logic_vector(to_unsigned( 95,8)),
			3525 => std_logic_vector(to_unsigned( 159,8)),
			3526 => std_logic_vector(to_unsigned( 12,8)),
			3527 => std_logic_vector(to_unsigned( 96,8)),
			3528 => std_logic_vector(to_unsigned( 133,8)),
			3529 => std_logic_vector(to_unsigned( 133,8)),
			3530 => std_logic_vector(to_unsigned( 133,8)),
			3531 => std_logic_vector(to_unsigned( 235,8)),
			3532 => std_logic_vector(to_unsigned( 45,8)),
			3533 => std_logic_vector(to_unsigned( 202,8)),
			3534 => std_logic_vector(to_unsigned( 168,8)),
			3535 => std_logic_vector(to_unsigned( 63,8)),
			3536 => std_logic_vector(to_unsigned( 234,8)),
			3537 => std_logic_vector(to_unsigned( 250,8)),
			3538 => std_logic_vector(to_unsigned( 254,8)),
			3539 => std_logic_vector(to_unsigned( 6,8)),
			3540 => std_logic_vector(to_unsigned( 117,8)),
			3541 => std_logic_vector(to_unsigned( 7,8)),
			3542 => std_logic_vector(to_unsigned( 57,8)),
			3543 => std_logic_vector(to_unsigned( 151,8)),
			3544 => std_logic_vector(to_unsigned( 135,8)),
			3545 => std_logic_vector(to_unsigned( 147,8)),
			3546 => std_logic_vector(to_unsigned( 137,8)),
			3547 => std_logic_vector(to_unsigned( 76,8)),
			3548 => std_logic_vector(to_unsigned( 75,8)),
			3549 => std_logic_vector(to_unsigned( 210,8)),
			3550 => std_logic_vector(to_unsigned( 234,8)),
			3551 => std_logic_vector(to_unsigned( 33,8)),
			3552 => std_logic_vector(to_unsigned( 150,8)),
			3553 => std_logic_vector(to_unsigned( 68,8)),
			3554 => std_logic_vector(to_unsigned( 76,8)),
			3555 => std_logic_vector(to_unsigned( 92,8)),
			3556 => std_logic_vector(to_unsigned( 146,8)),
			3557 => std_logic_vector(to_unsigned( 142,8)),
			3558 => std_logic_vector(to_unsigned( 195,8)),
			3559 => std_logic_vector(to_unsigned( 13,8)),
			3560 => std_logic_vector(to_unsigned( 184,8)),
			3561 => std_logic_vector(to_unsigned( 94,8)),
			3562 => std_logic_vector(to_unsigned( 121,8)),
			3563 => std_logic_vector(to_unsigned( 140,8)),
			3564 => std_logic_vector(to_unsigned( 249,8)),
			3565 => std_logic_vector(to_unsigned( 8,8)),
			3566 => std_logic_vector(to_unsigned( 94,8)),
			3567 => std_logic_vector(to_unsigned( 86,8)),
			3568 => std_logic_vector(to_unsigned( 239,8)),
			3569 => std_logic_vector(to_unsigned( 165,8)),
			3570 => std_logic_vector(to_unsigned( 254,8)),
			3571 => std_logic_vector(to_unsigned( 90,8)),
			3572 => std_logic_vector(to_unsigned( 14,8)),
			3573 => std_logic_vector(to_unsigned( 8,8)),
			3574 => std_logic_vector(to_unsigned( 84,8)),
			3575 => std_logic_vector(to_unsigned( 118,8)),
			3576 => std_logic_vector(to_unsigned( 143,8)),
			3577 => std_logic_vector(to_unsigned( 244,8)),
			3578 => std_logic_vector(to_unsigned( 173,8)),
			3579 => std_logic_vector(to_unsigned( 76,8)),
			3580 => std_logic_vector(to_unsigned( 137,8)),
			3581 => std_logic_vector(to_unsigned( 16,8)),
			3582 => std_logic_vector(to_unsigned( 47,8)),
			3583 => std_logic_vector(to_unsigned( 112,8)),
			3584 => std_logic_vector(to_unsigned( 117,8)),
			3585 => std_logic_vector(to_unsigned( 203,8)),
			3586 => std_logic_vector(to_unsigned( 105,8)),
			3587 => std_logic_vector(to_unsigned( 177,8)),
			3588 => std_logic_vector(to_unsigned( 4,8)),
			3589 => std_logic_vector(to_unsigned( 69,8)),
			3590 => std_logic_vector(to_unsigned( 181,8)),
			3591 => std_logic_vector(to_unsigned( 6,8)),
			3592 => std_logic_vector(to_unsigned( 95,8)),
			3593 => std_logic_vector(to_unsigned( 76,8)),
			3594 => std_logic_vector(to_unsigned( 185,8)),
			3595 => std_logic_vector(to_unsigned( 53,8)),
			3596 => std_logic_vector(to_unsigned( 41,8)),
			3597 => std_logic_vector(to_unsigned( 212,8)),
			3598 => std_logic_vector(to_unsigned( 111,8)),
			3599 => std_logic_vector(to_unsigned( 194,8)),
			3600 => std_logic_vector(to_unsigned( 80,8)),
			3601 => std_logic_vector(to_unsigned( 53,8)),
			3602 => std_logic_vector(to_unsigned( 114,8)),
			3603 => std_logic_vector(to_unsigned( 94,8)),
			3604 => std_logic_vector(to_unsigned( 174,8)),
			3605 => std_logic_vector(to_unsigned( 226,8)),
			3606 => std_logic_vector(to_unsigned( 33,8)),
			3607 => std_logic_vector(to_unsigned( 155,8)),
			3608 => std_logic_vector(to_unsigned( 124,8)),
			3609 => std_logic_vector(to_unsigned( 111,8)),
			3610 => std_logic_vector(to_unsigned( 117,8)),
			3611 => std_logic_vector(to_unsigned( 94,8)),
			3612 => std_logic_vector(to_unsigned( 216,8)),
			3613 => std_logic_vector(to_unsigned( 137,8)),
			3614 => std_logic_vector(to_unsigned( 81,8)),
			3615 => std_logic_vector(to_unsigned( 121,8)),
			3616 => std_logic_vector(to_unsigned( 17,8)),
			3617 => std_logic_vector(to_unsigned( 197,8)),
			3618 => std_logic_vector(to_unsigned( 15,8)),
			3619 => std_logic_vector(to_unsigned( 208,8)),
			3620 => std_logic_vector(to_unsigned( 104,8)),
			3621 => std_logic_vector(to_unsigned( 18,8)),
			3622 => std_logic_vector(to_unsigned( 63,8)),
			3623 => std_logic_vector(to_unsigned( 25,8)),
			3624 => std_logic_vector(to_unsigned( 188,8)),
			3625 => std_logic_vector(to_unsigned( 240,8)),
			3626 => std_logic_vector(to_unsigned( 92,8)),
			3627 => std_logic_vector(to_unsigned( 22,8)),
			3628 => std_logic_vector(to_unsigned( 223,8)),
			3629 => std_logic_vector(to_unsigned( 30,8)),
			3630 => std_logic_vector(to_unsigned( 119,8)),
			3631 => std_logic_vector(to_unsigned( 96,8)),
			3632 => std_logic_vector(to_unsigned( 174,8)),
			3633 => std_logic_vector(to_unsigned( 165,8)),
			3634 => std_logic_vector(to_unsigned( 253,8)),
			3635 => std_logic_vector(to_unsigned( 22,8)),
			3636 => std_logic_vector(to_unsigned( 79,8)),
			3637 => std_logic_vector(to_unsigned( 137,8)),
			3638 => std_logic_vector(to_unsigned( 153,8)),
			3639 => std_logic_vector(to_unsigned( 188,8)),
			3640 => std_logic_vector(to_unsigned( 55,8)),
			3641 => std_logic_vector(to_unsigned( 107,8)),
			3642 => std_logic_vector(to_unsigned( 235,8)),
			3643 => std_logic_vector(to_unsigned( 10,8)),
			3644 => std_logic_vector(to_unsigned( 251,8)),
			3645 => std_logic_vector(to_unsigned( 85,8)),
			3646 => std_logic_vector(to_unsigned( 220,8)),
			3647 => std_logic_vector(to_unsigned( 196,8)),
			3648 => std_logic_vector(to_unsigned( 204,8)),
			3649 => std_logic_vector(to_unsigned( 197,8)),
			3650 => std_logic_vector(to_unsigned( 247,8)),
			3651 => std_logic_vector(to_unsigned( 236,8)),
			3652 => std_logic_vector(to_unsigned( 137,8)),
			3653 => std_logic_vector(to_unsigned( 80,8)),
			3654 => std_logic_vector(to_unsigned( 184,8)),
			3655 => std_logic_vector(to_unsigned( 131,8)),
			3656 => std_logic_vector(to_unsigned( 33,8)),
			3657 => std_logic_vector(to_unsigned( 82,8)),
			3658 => std_logic_vector(to_unsigned( 184,8)),
			3659 => std_logic_vector(to_unsigned( 24,8)),
			3660 => std_logic_vector(to_unsigned( 180,8)),
			3661 => std_logic_vector(to_unsigned( 163,8)),
			3662 => std_logic_vector(to_unsigned( 47,8)),
			3663 => std_logic_vector(to_unsigned( 63,8)),
			3664 => std_logic_vector(to_unsigned( 33,8)),
			3665 => std_logic_vector(to_unsigned( 215,8)),
			3666 => std_logic_vector(to_unsigned( 25,8)),
			3667 => std_logic_vector(to_unsigned( 193,8)),
			3668 => std_logic_vector(to_unsigned( 48,8)),
			3669 => std_logic_vector(to_unsigned( 194,8)),
			3670 => std_logic_vector(to_unsigned( 106,8)),
			3671 => std_logic_vector(to_unsigned( 42,8)),
			3672 => std_logic_vector(to_unsigned( 124,8)),
			3673 => std_logic_vector(to_unsigned( 119,8)),
			3674 => std_logic_vector(to_unsigned( 187,8)),
			3675 => std_logic_vector(to_unsigned( 114,8)),
			3676 => std_logic_vector(to_unsigned( 230,8)),
			3677 => std_logic_vector(to_unsigned( 221,8)),
			3678 => std_logic_vector(to_unsigned( 85,8)),
			3679 => std_logic_vector(to_unsigned( 105,8)),
			3680 => std_logic_vector(to_unsigned( 8,8)),
			3681 => std_logic_vector(to_unsigned( 44,8)),
			3682 => std_logic_vector(to_unsigned( 192,8)),
			3683 => std_logic_vector(to_unsigned( 208,8)),
			3684 => std_logic_vector(to_unsigned( 15,8)),
			3685 => std_logic_vector(to_unsigned( 29,8)),
			3686 => std_logic_vector(to_unsigned( 88,8)),
			3687 => std_logic_vector(to_unsigned( 240,8)),
			3688 => std_logic_vector(to_unsigned( 30,8)),
			3689 => std_logic_vector(to_unsigned( 56,8)),
			3690 => std_logic_vector(to_unsigned( 11,8)),
			3691 => std_logic_vector(to_unsigned( 38,8)),
			3692 => std_logic_vector(to_unsigned( 202,8)),
			3693 => std_logic_vector(to_unsigned( 201,8)),
			3694 => std_logic_vector(to_unsigned( 226,8)),
			3695 => std_logic_vector(to_unsigned( 78,8)),
			3696 => std_logic_vector(to_unsigned( 30,8)),
			3697 => std_logic_vector(to_unsigned( 77,8)),
			3698 => std_logic_vector(to_unsigned( 126,8)),
			3699 => std_logic_vector(to_unsigned( 172,8)),
			3700 => std_logic_vector(to_unsigned( 185,8)),
			3701 => std_logic_vector(to_unsigned( 141,8)),
			3702 => std_logic_vector(to_unsigned( 116,8)),
			3703 => std_logic_vector(to_unsigned( 89,8)),
			3704 => std_logic_vector(to_unsigned( 89,8)),
			3705 => std_logic_vector(to_unsigned( 18,8)),
			3706 => std_logic_vector(to_unsigned( 93,8)),
			3707 => std_logic_vector(to_unsigned( 135,8)),
			3708 => std_logic_vector(to_unsigned( 121,8)),
			3709 => std_logic_vector(to_unsigned( 20,8)),
			3710 => std_logic_vector(to_unsigned( 197,8)),
			3711 => std_logic_vector(to_unsigned( 63,8)),
			3712 => std_logic_vector(to_unsigned( 3,8)),
			3713 => std_logic_vector(to_unsigned( 142,8)),
			3714 => std_logic_vector(to_unsigned( 131,8)),
			3715 => std_logic_vector(to_unsigned( 204,8)),
			3716 => std_logic_vector(to_unsigned( 229,8)),
			3717 => std_logic_vector(to_unsigned( 20,8)),
			3718 => std_logic_vector(to_unsigned( 13,8)),
			3719 => std_logic_vector(to_unsigned( 248,8)),
			3720 => std_logic_vector(to_unsigned( 1,8)),
			3721 => std_logic_vector(to_unsigned( 22,8)),
			3722 => std_logic_vector(to_unsigned( 66,8)),
			3723 => std_logic_vector(to_unsigned( 132,8)),
			3724 => std_logic_vector(to_unsigned( 193,8)),
			3725 => std_logic_vector(to_unsigned( 8,8)),
			3726 => std_logic_vector(to_unsigned( 64,8)),
			3727 => std_logic_vector(to_unsigned( 203,8)),
			3728 => std_logic_vector(to_unsigned( 172,8)),
			3729 => std_logic_vector(to_unsigned( 80,8)),
			3730 => std_logic_vector(to_unsigned( 43,8)),
			3731 => std_logic_vector(to_unsigned( 158,8)),
			3732 => std_logic_vector(to_unsigned( 106,8)),
			3733 => std_logic_vector(to_unsigned( 124,8)),
			3734 => std_logic_vector(to_unsigned( 155,8)),
			3735 => std_logic_vector(to_unsigned( 145,8)),
			3736 => std_logic_vector(to_unsigned( 159,8)),
			3737 => std_logic_vector(to_unsigned( 242,8)),
			3738 => std_logic_vector(to_unsigned( 122,8)),
			3739 => std_logic_vector(to_unsigned( 174,8)),
			3740 => std_logic_vector(to_unsigned( 25,8)),
			3741 => std_logic_vector(to_unsigned( 151,8)),
			3742 => std_logic_vector(to_unsigned( 35,8)),
			3743 => std_logic_vector(to_unsigned( 177,8)),
			3744 => std_logic_vector(to_unsigned( 20,8)),
			3745 => std_logic_vector(to_unsigned( 175,8)),
			3746 => std_logic_vector(to_unsigned( 55,8)),
			3747 => std_logic_vector(to_unsigned( 44,8)),
			3748 => std_logic_vector(to_unsigned( 57,8)),
			3749 => std_logic_vector(to_unsigned( 3,8)),
			3750 => std_logic_vector(to_unsigned( 170,8)),
			3751 => std_logic_vector(to_unsigned( 197,8)),
			3752 => std_logic_vector(to_unsigned( 152,8)),
			3753 => std_logic_vector(to_unsigned( 29,8)),
			3754 => std_logic_vector(to_unsigned( 150,8)),
			3755 => std_logic_vector(to_unsigned( 39,8)),
			3756 => std_logic_vector(to_unsigned( 13,8)),
			3757 => std_logic_vector(to_unsigned( 137,8)),
			3758 => std_logic_vector(to_unsigned( 177,8)),
			3759 => std_logic_vector(to_unsigned( 209,8)),
			3760 => std_logic_vector(to_unsigned( 226,8)),
			3761 => std_logic_vector(to_unsigned( 121,8)),
			3762 => std_logic_vector(to_unsigned( 134,8)),
			3763 => std_logic_vector(to_unsigned( 61,8)),
			3764 => std_logic_vector(to_unsigned( 85,8)),
			3765 => std_logic_vector(to_unsigned( 186,8)),
			3766 => std_logic_vector(to_unsigned( 177,8)),
			3767 => std_logic_vector(to_unsigned( 228,8)),
			3768 => std_logic_vector(to_unsigned( 55,8)),
			3769 => std_logic_vector(to_unsigned( 117,8)),
			3770 => std_logic_vector(to_unsigned( 18,8)),
			3771 => std_logic_vector(to_unsigned( 226,8)),
			3772 => std_logic_vector(to_unsigned( 46,8)),
			3773 => std_logic_vector(to_unsigned( 218,8)),
			3774 => std_logic_vector(to_unsigned( 253,8)),
			3775 => std_logic_vector(to_unsigned( 193,8)),
			3776 => std_logic_vector(to_unsigned( 85,8)),
			3777 => std_logic_vector(to_unsigned( 140,8)),
			3778 => std_logic_vector(to_unsigned( 220,8)),
			3779 => std_logic_vector(to_unsigned( 87,8)),
			3780 => std_logic_vector(to_unsigned( 140,8)),
			3781 => std_logic_vector(to_unsigned( 253,8)),
			3782 => std_logic_vector(to_unsigned( 79,8)),
			3783 => std_logic_vector(to_unsigned( 136,8)),
			3784 => std_logic_vector(to_unsigned( 78,8)),
			3785 => std_logic_vector(to_unsigned( 58,8)),
			3786 => std_logic_vector(to_unsigned( 31,8)),
			3787 => std_logic_vector(to_unsigned( 196,8)),
			3788 => std_logic_vector(to_unsigned( 215,8)),
			3789 => std_logic_vector(to_unsigned( 178,8)),
			3790 => std_logic_vector(to_unsigned( 156,8)),
			3791 => std_logic_vector(to_unsigned( 134,8)),
			3792 => std_logic_vector(to_unsigned( 90,8)),
			3793 => std_logic_vector(to_unsigned( 200,8)),
			3794 => std_logic_vector(to_unsigned( 121,8)),
			3795 => std_logic_vector(to_unsigned( 59,8)),
			3796 => std_logic_vector(to_unsigned( 58,8)),
			3797 => std_logic_vector(to_unsigned( 203,8)),
			3798 => std_logic_vector(to_unsigned( 66,8)),
			3799 => std_logic_vector(to_unsigned( 128,8)),
			3800 => std_logic_vector(to_unsigned( 222,8)),
			3801 => std_logic_vector(to_unsigned( 92,8)),
			3802 => std_logic_vector(to_unsigned( 130,8)),
			3803 => std_logic_vector(to_unsigned( 218,8)),
			3804 => std_logic_vector(to_unsigned( 0,8)),
			3805 => std_logic_vector(to_unsigned( 16,8)),
			3806 => std_logic_vector(to_unsigned( 17,8)),
			3807 => std_logic_vector(to_unsigned( 196,8)),
			3808 => std_logic_vector(to_unsigned( 177,8)),
			3809 => std_logic_vector(to_unsigned( 69,8)),
			3810 => std_logic_vector(to_unsigned( 213,8)),
			3811 => std_logic_vector(to_unsigned( 76,8)),
			3812 => std_logic_vector(to_unsigned( 5,8)),
			3813 => std_logic_vector(to_unsigned( 220,8)),
			3814 => std_logic_vector(to_unsigned( 89,8)),
			3815 => std_logic_vector(to_unsigned( 253,8)),
			3816 => std_logic_vector(to_unsigned( 107,8)),
			3817 => std_logic_vector(to_unsigned( 15,8)),
			3818 => std_logic_vector(to_unsigned( 3,8)),
			3819 => std_logic_vector(to_unsigned( 12,8)),
			3820 => std_logic_vector(to_unsigned( 173,8)),
			3821 => std_logic_vector(to_unsigned( 30,8)),
			3822 => std_logic_vector(to_unsigned( 170,8)),
			3823 => std_logic_vector(to_unsigned( 88,8)),
			3824 => std_logic_vector(to_unsigned( 150,8)),
			3825 => std_logic_vector(to_unsigned( 127,8)),
			3826 => std_logic_vector(to_unsigned( 64,8)),
			3827 => std_logic_vector(to_unsigned( 222,8)),
			3828 => std_logic_vector(to_unsigned( 247,8)),
			3829 => std_logic_vector(to_unsigned( 227,8)),
			3830 => std_logic_vector(to_unsigned( 174,8)),
			3831 => std_logic_vector(to_unsigned( 128,8)),
			3832 => std_logic_vector(to_unsigned( 118,8)),
			3833 => std_logic_vector(to_unsigned( 43,8)),
			3834 => std_logic_vector(to_unsigned( 91,8)),
			3835 => std_logic_vector(to_unsigned( 214,8)),
			3836 => std_logic_vector(to_unsigned( 171,8)),
			3837 => std_logic_vector(to_unsigned( 67,8)),
			3838 => std_logic_vector(to_unsigned( 43,8)),
			3839 => std_logic_vector(to_unsigned( 153,8)),
			3840 => std_logic_vector(to_unsigned( 113,8)),
			3841 => std_logic_vector(to_unsigned( 74,8)),
			3842 => std_logic_vector(to_unsigned( 132,8)),
			3843 => std_logic_vector(to_unsigned( 142,8)),
			3844 => std_logic_vector(to_unsigned( 47,8)),
			3845 => std_logic_vector(to_unsigned( 116,8)),
			3846 => std_logic_vector(to_unsigned( 34,8)),
			3847 => std_logic_vector(to_unsigned( 16,8)),
			3848 => std_logic_vector(to_unsigned( 25,8)),
			3849 => std_logic_vector(to_unsigned( 255,8)),
			3850 => std_logic_vector(to_unsigned( 168,8)),
			3851 => std_logic_vector(to_unsigned( 79,8)),
			3852 => std_logic_vector(to_unsigned( 181,8)),
			3853 => std_logic_vector(to_unsigned( 175,8)),
			3854 => std_logic_vector(to_unsigned( 99,8)),
			3855 => std_logic_vector(to_unsigned( 89,8)),
			3856 => std_logic_vector(to_unsigned( 13,8)),
			3857 => std_logic_vector(to_unsigned( 93,8)),
			3858 => std_logic_vector(to_unsigned( 171,8)),
			3859 => std_logic_vector(to_unsigned( 133,8)),
			3860 => std_logic_vector(to_unsigned( 101,8)),
			3861 => std_logic_vector(to_unsigned( 205,8)),
			3862 => std_logic_vector(to_unsigned( 176,8)),
			3863 => std_logic_vector(to_unsigned( 254,8)),
			3864 => std_logic_vector(to_unsigned( 61,8)),
			3865 => std_logic_vector(to_unsigned( 246,8)),
			3866 => std_logic_vector(to_unsigned( 181,8)),
			3867 => std_logic_vector(to_unsigned( 13,8)),
			3868 => std_logic_vector(to_unsigned( 229,8)),
			3869 => std_logic_vector(to_unsigned( 59,8)),
			3870 => std_logic_vector(to_unsigned( 113,8)),
			3871 => std_logic_vector(to_unsigned( 5,8)),
			3872 => std_logic_vector(to_unsigned( 16,8)),
			3873 => std_logic_vector(to_unsigned( 26,8)),
			3874 => std_logic_vector(to_unsigned( 200,8)),
			3875 => std_logic_vector(to_unsigned( 230,8)),
			3876 => std_logic_vector(to_unsigned( 145,8)),
			3877 => std_logic_vector(to_unsigned( 243,8)),
			3878 => std_logic_vector(to_unsigned( 8,8)),
			3879 => std_logic_vector(to_unsigned( 32,8)),
			3880 => std_logic_vector(to_unsigned( 215,8)),
			3881 => std_logic_vector(to_unsigned( 236,8)),
			3882 => std_logic_vector(to_unsigned( 96,8)),
			3883 => std_logic_vector(to_unsigned( 182,8)),
			3884 => std_logic_vector(to_unsigned( 82,8)),
			3885 => std_logic_vector(to_unsigned( 255,8)),
			3886 => std_logic_vector(to_unsigned( 110,8)),
			3887 => std_logic_vector(to_unsigned( 123,8)),
			3888 => std_logic_vector(to_unsigned( 69,8)),
			3889 => std_logic_vector(to_unsigned( 94,8)),
			3890 => std_logic_vector(to_unsigned( 22,8)),
			3891 => std_logic_vector(to_unsigned( 168,8)),
			3892 => std_logic_vector(to_unsigned( 28,8)),
			3893 => std_logic_vector(to_unsigned( 179,8)),
			3894 => std_logic_vector(to_unsigned( 157,8)),
			3895 => std_logic_vector(to_unsigned( 67,8)),
			3896 => std_logic_vector(to_unsigned( 55,8)),
			3897 => std_logic_vector(to_unsigned( 103,8)),
			3898 => std_logic_vector(to_unsigned( 70,8)),
			3899 => std_logic_vector(to_unsigned( 190,8)),
			3900 => std_logic_vector(to_unsigned( 164,8)),
			3901 => std_logic_vector(to_unsigned( 143,8)),
			3902 => std_logic_vector(to_unsigned( 219,8)),
			3903 => std_logic_vector(to_unsigned( 166,8)),
			3904 => std_logic_vector(to_unsigned( 118,8)),
			3905 => std_logic_vector(to_unsigned( 191,8)),
			3906 => std_logic_vector(to_unsigned( 150,8)),
			3907 => std_logic_vector(to_unsigned( 163,8)),
			3908 => std_logic_vector(to_unsigned( 36,8)),
			3909 => std_logic_vector(to_unsigned( 69,8)),
			3910 => std_logic_vector(to_unsigned( 173,8)),
			3911 => std_logic_vector(to_unsigned( 233,8)),
			3912 => std_logic_vector(to_unsigned( 234,8)),
			3913 => std_logic_vector(to_unsigned( 195,8)),
			3914 => std_logic_vector(to_unsigned( 88,8)),
			3915 => std_logic_vector(to_unsigned( 177,8)),
			3916 => std_logic_vector(to_unsigned( 206,8)),
			3917 => std_logic_vector(to_unsigned( 57,8)),
			3918 => std_logic_vector(to_unsigned( 185,8)),
			3919 => std_logic_vector(to_unsigned( 35,8)),
			3920 => std_logic_vector(to_unsigned( 23,8)),
			3921 => std_logic_vector(to_unsigned( 158,8)),
			3922 => std_logic_vector(to_unsigned( 20,8)),
			3923 => std_logic_vector(to_unsigned( 30,8)),
			3924 => std_logic_vector(to_unsigned( 35,8)),
			3925 => std_logic_vector(to_unsigned( 190,8)),
			3926 => std_logic_vector(to_unsigned( 61,8)),
			3927 => std_logic_vector(to_unsigned( 163,8)),
			3928 => std_logic_vector(to_unsigned( 204,8)),
			3929 => std_logic_vector(to_unsigned( 141,8)),
			3930 => std_logic_vector(to_unsigned( 134,8)),
			3931 => std_logic_vector(to_unsigned( 228,8)),
			3932 => std_logic_vector(to_unsigned( 231,8)),
			3933 => std_logic_vector(to_unsigned( 154,8)),
			3934 => std_logic_vector(to_unsigned( 241,8)),
			3935 => std_logic_vector(to_unsigned( 155,8)),
			3936 => std_logic_vector(to_unsigned( 112,8)),
			3937 => std_logic_vector(to_unsigned( 139,8)),
			3938 => std_logic_vector(to_unsigned( 127,8)),
			3939 => std_logic_vector(to_unsigned( 97,8)),
			3940 => std_logic_vector(to_unsigned( 197,8)),
			3941 => std_logic_vector(to_unsigned( 187,8)),
			3942 => std_logic_vector(to_unsigned( 234,8)),
			3943 => std_logic_vector(to_unsigned( 33,8)),
			3944 => std_logic_vector(to_unsigned( 20,8)),
			3945 => std_logic_vector(to_unsigned( 243,8)),
			3946 => std_logic_vector(to_unsigned( 254,8)),
			3947 => std_logic_vector(to_unsigned( 75,8)),
			3948 => std_logic_vector(to_unsigned( 200,8)),
			3949 => std_logic_vector(to_unsigned( 4,8)),
			3950 => std_logic_vector(to_unsigned( 207,8)),
			3951 => std_logic_vector(to_unsigned( 170,8)),
			3952 => std_logic_vector(to_unsigned( 35,8)),
			3953 => std_logic_vector(to_unsigned( 203,8)),
			3954 => std_logic_vector(to_unsigned( 119,8)),
			3955 => std_logic_vector(to_unsigned( 239,8)),
			3956 => std_logic_vector(to_unsigned( 135,8)),
			3957 => std_logic_vector(to_unsigned( 242,8)),
			3958 => std_logic_vector(to_unsigned( 10,8)),
			3959 => std_logic_vector(to_unsigned( 32,8)),
			3960 => std_logic_vector(to_unsigned( 134,8)),
			3961 => std_logic_vector(to_unsigned( 5,8)),
			3962 => std_logic_vector(to_unsigned( 145,8)),
			3963 => std_logic_vector(to_unsigned( 81,8)),
			3964 => std_logic_vector(to_unsigned( 116,8)),
			3965 => std_logic_vector(to_unsigned( 180,8)),
			3966 => std_logic_vector(to_unsigned( 36,8)),
			3967 => std_logic_vector(to_unsigned( 125,8)),
			3968 => std_logic_vector(to_unsigned( 48,8)),
			3969 => std_logic_vector(to_unsigned( 55,8)),
			3970 => std_logic_vector(to_unsigned( 199,8)),
			3971 => std_logic_vector(to_unsigned( 10,8)),
			3972 => std_logic_vector(to_unsigned( 238,8)),
			3973 => std_logic_vector(to_unsigned( 197,8)),
			3974 => std_logic_vector(to_unsigned( 196,8)),
			3975 => std_logic_vector(to_unsigned( 149,8)),
			3976 => std_logic_vector(to_unsigned( 99,8)),
			3977 => std_logic_vector(to_unsigned( 251,8)),
			3978 => std_logic_vector(to_unsigned( 30,8)),
			3979 => std_logic_vector(to_unsigned( 60,8)),
			3980 => std_logic_vector(to_unsigned( 122,8)),
			3981 => std_logic_vector(to_unsigned( 218,8)),
			3982 => std_logic_vector(to_unsigned( 40,8)),
			3983 => std_logic_vector(to_unsigned( 202,8)),
			3984 => std_logic_vector(to_unsigned( 60,8)),
			3985 => std_logic_vector(to_unsigned( 109,8)),
			3986 => std_logic_vector(to_unsigned( 74,8)),
			3987 => std_logic_vector(to_unsigned( 157,8)),
			3988 => std_logic_vector(to_unsigned( 234,8)),
			3989 => std_logic_vector(to_unsigned( 168,8)),
			3990 => std_logic_vector(to_unsigned( 1,8)),
			3991 => std_logic_vector(to_unsigned( 235,8)),
			3992 => std_logic_vector(to_unsigned( 102,8)),
			3993 => std_logic_vector(to_unsigned( 67,8)),
			3994 => std_logic_vector(to_unsigned( 165,8)),
			3995 => std_logic_vector(to_unsigned( 234,8)),
			3996 => std_logic_vector(to_unsigned( 137,8)),
			3997 => std_logic_vector(to_unsigned( 61,8)),
			3998 => std_logic_vector(to_unsigned( 33,8)),
			3999 => std_logic_vector(to_unsigned( 164,8)),
			4000 => std_logic_vector(to_unsigned( 11,8)),
			4001 => std_logic_vector(to_unsigned( 172,8)),
			4002 => std_logic_vector(to_unsigned( 131,8)),
			4003 => std_logic_vector(to_unsigned( 129,8)),
			4004 => std_logic_vector(to_unsigned( 78,8)),
			4005 => std_logic_vector(to_unsigned( 189,8)),
			4006 => std_logic_vector(to_unsigned( 146,8)),
			4007 => std_logic_vector(to_unsigned( 17,8)),
			4008 => std_logic_vector(to_unsigned( 103,8)),
			4009 => std_logic_vector(to_unsigned( 57,8)),
			4010 => std_logic_vector(to_unsigned( 237,8)),
			4011 => std_logic_vector(to_unsigned( 183,8)),
			4012 => std_logic_vector(to_unsigned( 142,8)),
			4013 => std_logic_vector(to_unsigned( 68,8)),
			4014 => std_logic_vector(to_unsigned( 5,8)),
			4015 => std_logic_vector(to_unsigned( 90,8)),
			4016 => std_logic_vector(to_unsigned( 89,8)),
			4017 => std_logic_vector(to_unsigned( 204,8)),
			4018 => std_logic_vector(to_unsigned( 159,8)),
			4019 => std_logic_vector(to_unsigned( 111,8)),
			4020 => std_logic_vector(to_unsigned( 117,8)),
			4021 => std_logic_vector(to_unsigned( 79,8)),
			4022 => std_logic_vector(to_unsigned( 203,8)),
			4023 => std_logic_vector(to_unsigned( 220,8)),
			4024 => std_logic_vector(to_unsigned( 120,8)),
			4025 => std_logic_vector(to_unsigned( 204,8)),
			4026 => std_logic_vector(to_unsigned( 252,8)),
			4027 => std_logic_vector(to_unsigned( 94,8)),
			4028 => std_logic_vector(to_unsigned( 161,8)),
			4029 => std_logic_vector(to_unsigned( 94,8)),
			4030 => std_logic_vector(to_unsigned( 23,8)),
			4031 => std_logic_vector(to_unsigned( 209,8)),
			4032 => std_logic_vector(to_unsigned( 120,8)),
			4033 => std_logic_vector(to_unsigned( 85,8)),
			4034 => std_logic_vector(to_unsigned( 6,8)),
			4035 => std_logic_vector(to_unsigned( 181,8)),
			4036 => std_logic_vector(to_unsigned( 139,8)),
			4037 => std_logic_vector(to_unsigned( 248,8)),
			4038 => std_logic_vector(to_unsigned( 125,8)),
			4039 => std_logic_vector(to_unsigned( 242,8)),
			4040 => std_logic_vector(to_unsigned( 146,8)),
			4041 => std_logic_vector(to_unsigned( 87,8)),
			4042 => std_logic_vector(to_unsigned( 111,8)),
			4043 => std_logic_vector(to_unsigned( 194,8)),
			4044 => std_logic_vector(to_unsigned( 232,8)),
			4045 => std_logic_vector(to_unsigned( 250,8)),
			4046 => std_logic_vector(to_unsigned( 110,8)),
			4047 => std_logic_vector(to_unsigned( 51,8)),
			4048 => std_logic_vector(to_unsigned( 146,8)),
			4049 => std_logic_vector(to_unsigned( 109,8)),
			4050 => std_logic_vector(to_unsigned( 182,8)),
			4051 => std_logic_vector(to_unsigned( 106,8)),
			4052 => std_logic_vector(to_unsigned( 214,8)),
			4053 => std_logic_vector(to_unsigned( 107,8)),
			4054 => std_logic_vector(to_unsigned( 239,8)),
			4055 => std_logic_vector(to_unsigned( 90,8)),
			4056 => std_logic_vector(to_unsigned( 119,8)),
			4057 => std_logic_vector(to_unsigned( 42,8)),
			4058 => std_logic_vector(to_unsigned( 224,8)),
			4059 => std_logic_vector(to_unsigned( 33,8)),
			4060 => std_logic_vector(to_unsigned( 252,8)),
			4061 => std_logic_vector(to_unsigned( 166,8)),
			4062 => std_logic_vector(to_unsigned( 111,8)),
			4063 => std_logic_vector(to_unsigned( 228,8)),
			4064 => std_logic_vector(to_unsigned( 96,8)),
			4065 => std_logic_vector(to_unsigned( 61,8)),
			4066 => std_logic_vector(to_unsigned( 23,8)),
			4067 => std_logic_vector(to_unsigned( 103,8)),
			4068 => std_logic_vector(to_unsigned( 21,8)),
			4069 => std_logic_vector(to_unsigned( 136,8)),
			4070 => std_logic_vector(to_unsigned( 1,8)),
			4071 => std_logic_vector(to_unsigned( 139,8)),
			4072 => std_logic_vector(to_unsigned( 229,8)),
			4073 => std_logic_vector(to_unsigned( 181,8)),
			4074 => std_logic_vector(to_unsigned( 195,8)),
			4075 => std_logic_vector(to_unsigned( 226,8)),
			4076 => std_logic_vector(to_unsigned( 122,8)),
			4077 => std_logic_vector(to_unsigned( 9,8)),
			4078 => std_logic_vector(to_unsigned( 10,8)),
			4079 => std_logic_vector(to_unsigned( 157,8)),
			4080 => std_logic_vector(to_unsigned( 57,8)),
			4081 => std_logic_vector(to_unsigned( 103,8)),
			4082 => std_logic_vector(to_unsigned( 202,8)),
			4083 => std_logic_vector(to_unsigned( 80,8)),
			4084 => std_logic_vector(to_unsigned( 185,8)),
			4085 => std_logic_vector(to_unsigned( 238,8)),
			4086 => std_logic_vector(to_unsigned( 231,8)),
			4087 => std_logic_vector(to_unsigned( 20,8)),
			4088 => std_logic_vector(to_unsigned( 218,8)),
			4089 => std_logic_vector(to_unsigned( 252,8)),
			4090 => std_logic_vector(to_unsigned( 36,8)),
			4091 => std_logic_vector(to_unsigned( 87,8)),
			4092 => std_logic_vector(to_unsigned( 72,8)),
			4093 => std_logic_vector(to_unsigned( 146,8)),
			4094 => std_logic_vector(to_unsigned( 63,8)),
			4095 => std_logic_vector(to_unsigned( 124,8)),
			4096 => std_logic_vector(to_unsigned( 199,8)),
			4097 => std_logic_vector(to_unsigned( 180,8)),
			4098 => std_logic_vector(to_unsigned( 212,8)),
			4099 => std_logic_vector(to_unsigned( 112,8)),
			4100 => std_logic_vector(to_unsigned( 73,8)),
			4101 => std_logic_vector(to_unsigned( 90,8)),
			4102 => std_logic_vector(to_unsigned( 146,8)),
			4103 => std_logic_vector(to_unsigned( 198,8)),
			4104 => std_logic_vector(to_unsigned( 167,8)),
			4105 => std_logic_vector(to_unsigned( 53,8)),
			4106 => std_logic_vector(to_unsigned( 223,8)),
			4107 => std_logic_vector(to_unsigned( 104,8)),
			4108 => std_logic_vector(to_unsigned( 250,8)),
			4109 => std_logic_vector(to_unsigned( 139,8)),
			4110 => std_logic_vector(to_unsigned( 119,8)),
			4111 => std_logic_vector(to_unsigned( 140,8)),
			4112 => std_logic_vector(to_unsigned( 194,8)),
			4113 => std_logic_vector(to_unsigned( 72,8)),
			4114 => std_logic_vector(to_unsigned( 91,8)),
			4115 => std_logic_vector(to_unsigned( 56,8)),
			4116 => std_logic_vector(to_unsigned( 105,8)),
			4117 => std_logic_vector(to_unsigned( 246,8)),
			4118 => std_logic_vector(to_unsigned( 76,8)),
			4119 => std_logic_vector(to_unsigned( 54,8)),
			4120 => std_logic_vector(to_unsigned( 233,8)),
			4121 => std_logic_vector(to_unsigned( 50,8)),
			4122 => std_logic_vector(to_unsigned( 221,8)),
			4123 => std_logic_vector(to_unsigned( 173,8)),
			4124 => std_logic_vector(to_unsigned( 122,8)),
			4125 => std_logic_vector(to_unsigned( 33,8)),
			4126 => std_logic_vector(to_unsigned( 69,8)),
			4127 => std_logic_vector(to_unsigned( 46,8)),
			4128 => std_logic_vector(to_unsigned( 241,8)),
			4129 => std_logic_vector(to_unsigned( 24,8)),
			4130 => std_logic_vector(to_unsigned( 157,8)),
			4131 => std_logic_vector(to_unsigned( 233,8)),
			4132 => std_logic_vector(to_unsigned( 84,8)),
			4133 => std_logic_vector(to_unsigned( 61,8)),
			4134 => std_logic_vector(to_unsigned( 88,8)),
			4135 => std_logic_vector(to_unsigned( 118,8)),
			4136 => std_logic_vector(to_unsigned( 63,8)),
			4137 => std_logic_vector(to_unsigned( 173,8)),
			4138 => std_logic_vector(to_unsigned( 175,8)),
			4139 => std_logic_vector(to_unsigned( 5,8)),
			4140 => std_logic_vector(to_unsigned( 110,8)),
			4141 => std_logic_vector(to_unsigned( 73,8)),
			4142 => std_logic_vector(to_unsigned( 45,8)),
			4143 => std_logic_vector(to_unsigned( 193,8)),
			4144 => std_logic_vector(to_unsigned( 222,8)),
			4145 => std_logic_vector(to_unsigned( 13,8)),
			4146 => std_logic_vector(to_unsigned( 122,8)),
			4147 => std_logic_vector(to_unsigned( 33,8)),
			4148 => std_logic_vector(to_unsigned( 29,8)),
			4149 => std_logic_vector(to_unsigned( 123,8)),
			4150 => std_logic_vector(to_unsigned( 20,8)),
			4151 => std_logic_vector(to_unsigned( 123,8)),
			4152 => std_logic_vector(to_unsigned( 50,8)),
			4153 => std_logic_vector(to_unsigned( 37,8)),
			4154 => std_logic_vector(to_unsigned( 251,8)),
			4155 => std_logic_vector(to_unsigned( 86,8)),
			4156 => std_logic_vector(to_unsigned( 230,8)),
			4157 => std_logic_vector(to_unsigned( 232,8)),
			4158 => std_logic_vector(to_unsigned( 186,8)),
			4159 => std_logic_vector(to_unsigned( 78,8)),
			4160 => std_logic_vector(to_unsigned( 114,8)),
			4161 => std_logic_vector(to_unsigned( 160,8)),
			4162 => std_logic_vector(to_unsigned( 9,8)),
			4163 => std_logic_vector(to_unsigned( 29,8)),
			4164 => std_logic_vector(to_unsigned( 234,8)),
			4165 => std_logic_vector(to_unsigned( 110,8)),
			4166 => std_logic_vector(to_unsigned( 23,8)),
			4167 => std_logic_vector(to_unsigned( 200,8)),
			4168 => std_logic_vector(to_unsigned( 183,8)),
			4169 => std_logic_vector(to_unsigned( 96,8)),
			4170 => std_logic_vector(to_unsigned( 26,8)),
			4171 => std_logic_vector(to_unsigned( 43,8)),
			4172 => std_logic_vector(to_unsigned( 53,8)),
			4173 => std_logic_vector(to_unsigned( 210,8)),
			4174 => std_logic_vector(to_unsigned( 203,8)),
			4175 => std_logic_vector(to_unsigned( 71,8)),
			4176 => std_logic_vector(to_unsigned( 205,8)),
			4177 => std_logic_vector(to_unsigned( 218,8)),
			4178 => std_logic_vector(to_unsigned( 182,8)),
			4179 => std_logic_vector(to_unsigned( 249,8)),
			4180 => std_logic_vector(to_unsigned( 219,8)),
			4181 => std_logic_vector(to_unsigned( 43,8)),
			4182 => std_logic_vector(to_unsigned( 187,8)),
			4183 => std_logic_vector(to_unsigned( 37,8)),
			4184 => std_logic_vector(to_unsigned( 250,8)),
			4185 => std_logic_vector(to_unsigned( 149,8)),
			4186 => std_logic_vector(to_unsigned( 241,8)),
			4187 => std_logic_vector(to_unsigned( 80,8)),
			4188 => std_logic_vector(to_unsigned( 94,8)),
			4189 => std_logic_vector(to_unsigned( 19,8)),
			4190 => std_logic_vector(to_unsigned( 120,8)),
			4191 => std_logic_vector(to_unsigned( 155,8)),
			4192 => std_logic_vector(to_unsigned( 131,8)),
			4193 => std_logic_vector(to_unsigned( 40,8)),
			4194 => std_logic_vector(to_unsigned( 40,8)),
			4195 => std_logic_vector(to_unsigned( 124,8)),
			4196 => std_logic_vector(to_unsigned( 53,8)),
			4197 => std_logic_vector(to_unsigned( 92,8)),
			4198 => std_logic_vector(to_unsigned( 225,8)),
			4199 => std_logic_vector(to_unsigned( 191,8)),
			4200 => std_logic_vector(to_unsigned( 233,8)),
			4201 => std_logic_vector(to_unsigned( 252,8)),
			4202 => std_logic_vector(to_unsigned( 34,8)),
			4203 => std_logic_vector(to_unsigned( 167,8)),
			4204 => std_logic_vector(to_unsigned( 211,8)),
			4205 => std_logic_vector(to_unsigned( 5,8)),
			4206 => std_logic_vector(to_unsigned( 195,8)),
			4207 => std_logic_vector(to_unsigned( 178,8)),
			4208 => std_logic_vector(to_unsigned( 67,8)),
			4209 => std_logic_vector(to_unsigned( 244,8)),
			4210 => std_logic_vector(to_unsigned( 139,8)),
			4211 => std_logic_vector(to_unsigned( 209,8)),
			4212 => std_logic_vector(to_unsigned( 74,8)),
			4213 => std_logic_vector(to_unsigned( 9,8)),
			4214 => std_logic_vector(to_unsigned( 29,8)),
			4215 => std_logic_vector(to_unsigned( 147,8)),
			4216 => std_logic_vector(to_unsigned( 26,8)),
			4217 => std_logic_vector(to_unsigned( 181,8)),
			4218 => std_logic_vector(to_unsigned( 170,8)),
			4219 => std_logic_vector(to_unsigned( 127,8)),
			4220 => std_logic_vector(to_unsigned( 193,8)),
			4221 => std_logic_vector(to_unsigned( 151,8)),
			4222 => std_logic_vector(to_unsigned( 65,8)),
			4223 => std_logic_vector(to_unsigned( 211,8)),
			4224 => std_logic_vector(to_unsigned( 136,8)),
			4225 => std_logic_vector(to_unsigned( 80,8)),
			4226 => std_logic_vector(to_unsigned( 232,8)),
			4227 => std_logic_vector(to_unsigned( 172,8)),
			4228 => std_logic_vector(to_unsigned( 142,8)),
			4229 => std_logic_vector(to_unsigned( 58,8)),
			4230 => std_logic_vector(to_unsigned( 225,8)),
			4231 => std_logic_vector(to_unsigned( 25,8)),
			4232 => std_logic_vector(to_unsigned( 188,8)),
			4233 => std_logic_vector(to_unsigned( 249,8)),
			4234 => std_logic_vector(to_unsigned( 73,8)),
			4235 => std_logic_vector(to_unsigned( 56,8)),
			4236 => std_logic_vector(to_unsigned( 34,8)),
			4237 => std_logic_vector(to_unsigned( 112,8)),
			4238 => std_logic_vector(to_unsigned( 106,8)),
			4239 => std_logic_vector(to_unsigned( 17,8)),
			4240 => std_logic_vector(to_unsigned( 126,8)),
			4241 => std_logic_vector(to_unsigned( 217,8)),
			4242 => std_logic_vector(to_unsigned( 153,8)),
			4243 => std_logic_vector(to_unsigned( 25,8)),
			4244 => std_logic_vector(to_unsigned( 169,8)),
			4245 => std_logic_vector(to_unsigned( 90,8)),
			4246 => std_logic_vector(to_unsigned( 253,8)),
			4247 => std_logic_vector(to_unsigned( 29,8)),
			4248 => std_logic_vector(to_unsigned( 87,8)),
			4249 => std_logic_vector(to_unsigned( 251,8)),
			4250 => std_logic_vector(to_unsigned( 164,8)),
			4251 => std_logic_vector(to_unsigned( 251,8)),
			4252 => std_logic_vector(to_unsigned( 146,8)),
			4253 => std_logic_vector(to_unsigned( 201,8)),
			4254 => std_logic_vector(to_unsigned( 92,8)),
			4255 => std_logic_vector(to_unsigned( 101,8)),
			4256 => std_logic_vector(to_unsigned( 234,8)),
			4257 => std_logic_vector(to_unsigned( 110,8)),
			4258 => std_logic_vector(to_unsigned( 12,8)),
			4259 => std_logic_vector(to_unsigned( 9,8)),
			4260 => std_logic_vector(to_unsigned( 76,8)),
			4261 => std_logic_vector(to_unsigned( 173,8)),
			4262 => std_logic_vector(to_unsigned( 242,8)),
			4263 => std_logic_vector(to_unsigned( 113,8)),
			4264 => std_logic_vector(to_unsigned( 106,8)),
			4265 => std_logic_vector(to_unsigned( 248,8)),
			4266 => std_logic_vector(to_unsigned( 105,8)),
			4267 => std_logic_vector(to_unsigned( 223,8)),
			4268 => std_logic_vector(to_unsigned( 46,8)),
			4269 => std_logic_vector(to_unsigned( 127,8)),
			4270 => std_logic_vector(to_unsigned( 60,8)),
			4271 => std_logic_vector(to_unsigned( 145,8)),
			4272 => std_logic_vector(to_unsigned( 109,8)),
			4273 => std_logic_vector(to_unsigned( 95,8)),
			4274 => std_logic_vector(to_unsigned( 6,8)),
			4275 => std_logic_vector(to_unsigned( 178,8)),
			4276 => std_logic_vector(to_unsigned( 244,8)),
			4277 => std_logic_vector(to_unsigned( 247,8)),
			4278 => std_logic_vector(to_unsigned( 218,8)),
			4279 => std_logic_vector(to_unsigned( 160,8)),
			4280 => std_logic_vector(to_unsigned( 89,8)),
			4281 => std_logic_vector(to_unsigned( 243,8)),
			4282 => std_logic_vector(to_unsigned( 183,8)),
			4283 => std_logic_vector(to_unsigned( 61,8)),
			4284 => std_logic_vector(to_unsigned( 232,8)),
			4285 => std_logic_vector(to_unsigned( 70,8)),
			4286 => std_logic_vector(to_unsigned( 34,8)),
			4287 => std_logic_vector(to_unsigned( 76,8)),
			4288 => std_logic_vector(to_unsigned( 85,8)),
			4289 => std_logic_vector(to_unsigned( 88,8)),
			4290 => std_logic_vector(to_unsigned( 62,8)),
			4291 => std_logic_vector(to_unsigned( 166,8)),
			4292 => std_logic_vector(to_unsigned( 67,8)),
			4293 => std_logic_vector(to_unsigned( 22,8)),
			4294 => std_logic_vector(to_unsigned( 101,8)),
			4295 => std_logic_vector(to_unsigned( 131,8)),
			4296 => std_logic_vector(to_unsigned( 191,8)),
			4297 => std_logic_vector(to_unsigned( 78,8)),
			4298 => std_logic_vector(to_unsigned( 227,8)),
			4299 => std_logic_vector(to_unsigned( 105,8)),
			4300 => std_logic_vector(to_unsigned( 130,8)),
			4301 => std_logic_vector(to_unsigned( 22,8)),
			4302 => std_logic_vector(to_unsigned( 194,8)),
			4303 => std_logic_vector(to_unsigned( 120,8)),
			4304 => std_logic_vector(to_unsigned( 99,8)),
			4305 => std_logic_vector(to_unsigned( 22,8)),
			4306 => std_logic_vector(to_unsigned( 254,8)),
			4307 => std_logic_vector(to_unsigned( 207,8)),
			4308 => std_logic_vector(to_unsigned( 70,8)),
			4309 => std_logic_vector(to_unsigned( 111,8)),
			4310 => std_logic_vector(to_unsigned( 195,8)),
			4311 => std_logic_vector(to_unsigned( 45,8)),
			4312 => std_logic_vector(to_unsigned( 177,8)),
			4313 => std_logic_vector(to_unsigned( 18,8)),
			4314 => std_logic_vector(to_unsigned( 203,8)),
			4315 => std_logic_vector(to_unsigned( 38,8)),
			4316 => std_logic_vector(to_unsigned( 14,8)),
			4317 => std_logic_vector(to_unsigned( 128,8)),
			4318 => std_logic_vector(to_unsigned( 80,8)),
			4319 => std_logic_vector(to_unsigned( 66,8)),
			4320 => std_logic_vector(to_unsigned( 99,8)),
			4321 => std_logic_vector(to_unsigned( 135,8)),
			4322 => std_logic_vector(to_unsigned( 55,8)),
			4323 => std_logic_vector(to_unsigned( 112,8)),
			4324 => std_logic_vector(to_unsigned( 168,8)),
			4325 => std_logic_vector(to_unsigned( 117,8)),
			4326 => std_logic_vector(to_unsigned( 6,8)),
			4327 => std_logic_vector(to_unsigned( 95,8)),
			4328 => std_logic_vector(to_unsigned( 139,8)),
			4329 => std_logic_vector(to_unsigned( 240,8)),
			4330 => std_logic_vector(to_unsigned( 75,8)),
			4331 => std_logic_vector(to_unsigned( 226,8)),
			4332 => std_logic_vector(to_unsigned( 123,8)),
			4333 => std_logic_vector(to_unsigned( 79,8)),
			4334 => std_logic_vector(to_unsigned( 84,8)),
			4335 => std_logic_vector(to_unsigned( 218,8)),
			4336 => std_logic_vector(to_unsigned( 58,8)),
			4337 => std_logic_vector(to_unsigned( 250,8)),
			4338 => std_logic_vector(to_unsigned( 107,8)),
			4339 => std_logic_vector(to_unsigned( 227,8)),
			4340 => std_logic_vector(to_unsigned( 31,8)),
			4341 => std_logic_vector(to_unsigned( 102,8)),
			4342 => std_logic_vector(to_unsigned( 191,8)),
			4343 => std_logic_vector(to_unsigned( 33,8)),
			4344 => std_logic_vector(to_unsigned( 168,8)),
			4345 => std_logic_vector(to_unsigned( 156,8)),
			4346 => std_logic_vector(to_unsigned( 135,8)),
			4347 => std_logic_vector(to_unsigned( 240,8)),
			4348 => std_logic_vector(to_unsigned( 58,8)),
			4349 => std_logic_vector(to_unsigned( 96,8)),
			4350 => std_logic_vector(to_unsigned( 57,8)),
			4351 => std_logic_vector(to_unsigned( 186,8)),
			4352 => std_logic_vector(to_unsigned( 184,8)),
			4353 => std_logic_vector(to_unsigned( 143,8)),
			4354 => std_logic_vector(to_unsigned( 207,8)),
			4355 => std_logic_vector(to_unsigned( 219,8)),
			4356 => std_logic_vector(to_unsigned( 140,8)),
			4357 => std_logic_vector(to_unsigned( 133,8)),
			4358 => std_logic_vector(to_unsigned( 175,8)),
			4359 => std_logic_vector(to_unsigned( 224,8)),
			4360 => std_logic_vector(to_unsigned( 72,8)),
			4361 => std_logic_vector(to_unsigned( 54,8)),
			4362 => std_logic_vector(to_unsigned( 191,8)),
			4363 => std_logic_vector(to_unsigned( 148,8)),
			4364 => std_logic_vector(to_unsigned( 8,8)),
			4365 => std_logic_vector(to_unsigned( 89,8)),
			4366 => std_logic_vector(to_unsigned( 57,8)),
			4367 => std_logic_vector(to_unsigned( 132,8)),
			4368 => std_logic_vector(to_unsigned( 235,8)),
			4369 => std_logic_vector(to_unsigned( 161,8)),
			4370 => std_logic_vector(to_unsigned( 98,8)),
			4371 => std_logic_vector(to_unsigned( 219,8)),
			4372 => std_logic_vector(to_unsigned( 28,8)),
			4373 => std_logic_vector(to_unsigned( 35,8)),
			4374 => std_logic_vector(to_unsigned( 172,8)),
			4375 => std_logic_vector(to_unsigned( 65,8)),
			4376 => std_logic_vector(to_unsigned( 64,8)),
			4377 => std_logic_vector(to_unsigned( 70,8)),
			4378 => std_logic_vector(to_unsigned( 234,8)),
			4379 => std_logic_vector(to_unsigned( 176,8)),
			4380 => std_logic_vector(to_unsigned( 68,8)),
			4381 => std_logic_vector(to_unsigned( 245,8)),
			4382 => std_logic_vector(to_unsigned( 200,8)),
			4383 => std_logic_vector(to_unsigned( 81,8)),
			4384 => std_logic_vector(to_unsigned( 157,8)),
			4385 => std_logic_vector(to_unsigned( 107,8)),
			4386 => std_logic_vector(to_unsigned( 191,8)),
			4387 => std_logic_vector(to_unsigned( 142,8)),
			4388 => std_logic_vector(to_unsigned( 3,8)),
			4389 => std_logic_vector(to_unsigned( 223,8)),
			4390 => std_logic_vector(to_unsigned( 84,8)),
			4391 => std_logic_vector(to_unsigned( 139,8)),
			4392 => std_logic_vector(to_unsigned( 10,8)),
			4393 => std_logic_vector(to_unsigned( 211,8)),
			4394 => std_logic_vector(to_unsigned( 113,8)),
			4395 => std_logic_vector(to_unsigned( 82,8)),
			4396 => std_logic_vector(to_unsigned( 44,8)),
			4397 => std_logic_vector(to_unsigned( 196,8)),
			4398 => std_logic_vector(to_unsigned( 176,8)),
			4399 => std_logic_vector(to_unsigned( 46,8)),
			4400 => std_logic_vector(to_unsigned( 15,8)),
			4401 => std_logic_vector(to_unsigned( 219,8)),
			4402 => std_logic_vector(to_unsigned( 154,8)),
			4403 => std_logic_vector(to_unsigned( 232,8)),
			4404 => std_logic_vector(to_unsigned( 187,8)),
			4405 => std_logic_vector(to_unsigned( 89,8)),
			4406 => std_logic_vector(to_unsigned( 180,8)),
			4407 => std_logic_vector(to_unsigned( 77,8)),
			4408 => std_logic_vector(to_unsigned( 184,8)),
			4409 => std_logic_vector(to_unsigned( 5,8)),
			4410 => std_logic_vector(to_unsigned( 113,8)),
			4411 => std_logic_vector(to_unsigned( 20,8)),
			4412 => std_logic_vector(to_unsigned( 79,8)),
			4413 => std_logic_vector(to_unsigned( 251,8)),
			4414 => std_logic_vector(to_unsigned( 1,8)),
			4415 => std_logic_vector(to_unsigned( 212,8)),
			4416 => std_logic_vector(to_unsigned( 197,8)),
			4417 => std_logic_vector(to_unsigned( 165,8)),
			4418 => std_logic_vector(to_unsigned( 105,8)),
			4419 => std_logic_vector(to_unsigned( 179,8)),
			4420 => std_logic_vector(to_unsigned( 156,8)),
			4421 => std_logic_vector(to_unsigned( 89,8)),
			4422 => std_logic_vector(to_unsigned( 135,8)),
			4423 => std_logic_vector(to_unsigned( 213,8)),
			4424 => std_logic_vector(to_unsigned( 211,8)),
			4425 => std_logic_vector(to_unsigned( 111,8)),
			4426 => std_logic_vector(to_unsigned( 68,8)),
			4427 => std_logic_vector(to_unsigned( 158,8)),
			4428 => std_logic_vector(to_unsigned( 117,8)),
			4429 => std_logic_vector(to_unsigned( 89,8)),
			4430 => std_logic_vector(to_unsigned( 68,8)),
			4431 => std_logic_vector(to_unsigned( 122,8)),
			4432 => std_logic_vector(to_unsigned( 155,8)),
			4433 => std_logic_vector(to_unsigned( 51,8)),
			4434 => std_logic_vector(to_unsigned( 220,8)),
			4435 => std_logic_vector(to_unsigned( 158,8)),
			4436 => std_logic_vector(to_unsigned( 106,8)),
			4437 => std_logic_vector(to_unsigned( 19,8)),
			4438 => std_logic_vector(to_unsigned( 69,8)),
			4439 => std_logic_vector(to_unsigned( 217,8)),
			4440 => std_logic_vector(to_unsigned( 251,8)),
			4441 => std_logic_vector(to_unsigned( 98,8)),
			4442 => std_logic_vector(to_unsigned( 155,8)),
			4443 => std_logic_vector(to_unsigned( 209,8)),
			4444 => std_logic_vector(to_unsigned( 121,8)),
			4445 => std_logic_vector(to_unsigned( 141,8)),
			4446 => std_logic_vector(to_unsigned( 146,8)),
			4447 => std_logic_vector(to_unsigned( 154,8)),
			4448 => std_logic_vector(to_unsigned( 3,8)),
			4449 => std_logic_vector(to_unsigned( 80,8)),
			4450 => std_logic_vector(to_unsigned( 202,8)),
			4451 => std_logic_vector(to_unsigned( 217,8)),
			4452 => std_logic_vector(to_unsigned( 229,8)),
			4453 => std_logic_vector(to_unsigned( 244,8)),
			4454 => std_logic_vector(to_unsigned( 186,8)),
			4455 => std_logic_vector(to_unsigned( 72,8)),
			4456 => std_logic_vector(to_unsigned( 131,8)),
			4457 => std_logic_vector(to_unsigned( 223,8)),
			4458 => std_logic_vector(to_unsigned( 156,8)),
			4459 => std_logic_vector(to_unsigned( 63,8)),
			4460 => std_logic_vector(to_unsigned( 101,8)),
			4461 => std_logic_vector(to_unsigned( 50,8)),
			4462 => std_logic_vector(to_unsigned( 202,8)),
			4463 => std_logic_vector(to_unsigned( 202,8)),
			4464 => std_logic_vector(to_unsigned( 191,8)),
			4465 => std_logic_vector(to_unsigned( 230,8)),
			4466 => std_logic_vector(to_unsigned( 168,8)),
			4467 => std_logic_vector(to_unsigned( 54,8)),
			4468 => std_logic_vector(to_unsigned( 178,8)),
			4469 => std_logic_vector(to_unsigned( 181,8)),
			4470 => std_logic_vector(to_unsigned( 23,8)),
			4471 => std_logic_vector(to_unsigned( 197,8)),
			4472 => std_logic_vector(to_unsigned( 185,8)),
			4473 => std_logic_vector(to_unsigned( 81,8)),
			4474 => std_logic_vector(to_unsigned( 255,8)),
			4475 => std_logic_vector(to_unsigned( 111,8)),
			4476 => std_logic_vector(to_unsigned( 230,8)),
			4477 => std_logic_vector(to_unsigned( 102,8)),
			4478 => std_logic_vector(to_unsigned( 54,8)),
			4479 => std_logic_vector(to_unsigned( 214,8)),
			4480 => std_logic_vector(to_unsigned( 177,8)),
			4481 => std_logic_vector(to_unsigned( 215,8)),
			4482 => std_logic_vector(to_unsigned( 122,8)),
			4483 => std_logic_vector(to_unsigned( 92,8)),
			4484 => std_logic_vector(to_unsigned( 123,8)),
			4485 => std_logic_vector(to_unsigned( 7,8)),
			4486 => std_logic_vector(to_unsigned( 84,8)),
			4487 => std_logic_vector(to_unsigned( 171,8)),
			4488 => std_logic_vector(to_unsigned( 251,8)),
			4489 => std_logic_vector(to_unsigned( 78,8)),
			4490 => std_logic_vector(to_unsigned( 175,8)),
			4491 => std_logic_vector(to_unsigned( 115,8)),
			4492 => std_logic_vector(to_unsigned( 183,8)),
			4493 => std_logic_vector(to_unsigned( 36,8)),
			4494 => std_logic_vector(to_unsigned( 51,8)),
			4495 => std_logic_vector(to_unsigned( 212,8)),
			4496 => std_logic_vector(to_unsigned( 116,8)),
			4497 => std_logic_vector(to_unsigned( 230,8)),
			4498 => std_logic_vector(to_unsigned( 202,8)),
			4499 => std_logic_vector(to_unsigned( 110,8)),
			4500 => std_logic_vector(to_unsigned( 230,8)),
			4501 => std_logic_vector(to_unsigned( 80,8)),
			4502 => std_logic_vector(to_unsigned( 71,8)),
			4503 => std_logic_vector(to_unsigned( 142,8)),
			4504 => std_logic_vector(to_unsigned( 20,8)),
			4505 => std_logic_vector(to_unsigned( 5,8)),
			4506 => std_logic_vector(to_unsigned( 113,8)),
			4507 => std_logic_vector(to_unsigned( 164,8)),
			4508 => std_logic_vector(to_unsigned( 243,8)),
			4509 => std_logic_vector(to_unsigned( 233,8)),
			4510 => std_logic_vector(to_unsigned( 214,8)),
			4511 => std_logic_vector(to_unsigned( 197,8)),
			4512 => std_logic_vector(to_unsigned( 103,8)),
			4513 => std_logic_vector(to_unsigned( 226,8)),
			4514 => std_logic_vector(to_unsigned( 99,8)),
			4515 => std_logic_vector(to_unsigned( 248,8)),
			4516 => std_logic_vector(to_unsigned( 209,8)),
			4517 => std_logic_vector(to_unsigned( 98,8)),
			4518 => std_logic_vector(to_unsigned( 51,8)),
			4519 => std_logic_vector(to_unsigned( 132,8)),
			4520 => std_logic_vector(to_unsigned( 32,8)),
			4521 => std_logic_vector(to_unsigned( 197,8)),
			4522 => std_logic_vector(to_unsigned( 60,8)),
			4523 => std_logic_vector(to_unsigned( 21,8)),
			4524 => std_logic_vector(to_unsigned( 193,8)),
			4525 => std_logic_vector(to_unsigned( 55,8)),
			4526 => std_logic_vector(to_unsigned( 247,8)),
			4527 => std_logic_vector(to_unsigned( 161,8)),
			4528 => std_logic_vector(to_unsigned( 193,8)),
			4529 => std_logic_vector(to_unsigned( 35,8)),
			4530 => std_logic_vector(to_unsigned( 63,8)),
			4531 => std_logic_vector(to_unsigned( 194,8)),
			4532 => std_logic_vector(to_unsigned( 63,8)),
			4533 => std_logic_vector(to_unsigned( 152,8)),
			4534 => std_logic_vector(to_unsigned( 209,8)),
			4535 => std_logic_vector(to_unsigned( 20,8)),
			4536 => std_logic_vector(to_unsigned( 165,8)),
			4537 => std_logic_vector(to_unsigned( 145,8)),
			4538 => std_logic_vector(to_unsigned( 50,8)),
			4539 => std_logic_vector(to_unsigned( 26,8)),
			4540 => std_logic_vector(to_unsigned( 90,8)),
			4541 => std_logic_vector(to_unsigned( 170,8)),
			4542 => std_logic_vector(to_unsigned( 19,8)),
			4543 => std_logic_vector(to_unsigned( 223,8)),
			4544 => std_logic_vector(to_unsigned( 170,8)),
			4545 => std_logic_vector(to_unsigned( 100,8)),
			4546 => std_logic_vector(to_unsigned( 58,8)),
			4547 => std_logic_vector(to_unsigned( 203,8)),
			4548 => std_logic_vector(to_unsigned( 39,8)),
			4549 => std_logic_vector(to_unsigned( 215,8)),
			4550 => std_logic_vector(to_unsigned( 8,8)),
			4551 => std_logic_vector(to_unsigned( 180,8)),
			4552 => std_logic_vector(to_unsigned( 4,8)),
			4553 => std_logic_vector(to_unsigned( 184,8)),
			4554 => std_logic_vector(to_unsigned( 219,8)),
			4555 => std_logic_vector(to_unsigned( 235,8)),
			4556 => std_logic_vector(to_unsigned( 146,8)),
			4557 => std_logic_vector(to_unsigned( 93,8)),
			4558 => std_logic_vector(to_unsigned( 87,8)),
			4559 => std_logic_vector(to_unsigned( 166,8)),
			4560 => std_logic_vector(to_unsigned( 145,8)),
			4561 => std_logic_vector(to_unsigned( 215,8)),
			4562 => std_logic_vector(to_unsigned( 255,8)),
			4563 => std_logic_vector(to_unsigned( 155,8)),
			4564 => std_logic_vector(to_unsigned( 91,8)),
			4565 => std_logic_vector(to_unsigned( 10,8)),
			4566 => std_logic_vector(to_unsigned( 31,8)),
			4567 => std_logic_vector(to_unsigned( 151,8)),
			4568 => std_logic_vector(to_unsigned( 91,8)),
			4569 => std_logic_vector(to_unsigned( 176,8)),
			4570 => std_logic_vector(to_unsigned( 72,8)),
			4571 => std_logic_vector(to_unsigned( 128,8)),
			4572 => std_logic_vector(to_unsigned( 116,8)),
			4573 => std_logic_vector(to_unsigned( 195,8)),
			4574 => std_logic_vector(to_unsigned( 83,8)),
			4575 => std_logic_vector(to_unsigned( 196,8)),
			4576 => std_logic_vector(to_unsigned( 62,8)),
			4577 => std_logic_vector(to_unsigned( 190,8)),
			4578 => std_logic_vector(to_unsigned( 240,8)),
			4579 => std_logic_vector(to_unsigned( 213,8)),
			4580 => std_logic_vector(to_unsigned( 161,8)),
			4581 => std_logic_vector(to_unsigned( 89,8)),
			4582 => std_logic_vector(to_unsigned( 161,8)),
			4583 => std_logic_vector(to_unsigned( 163,8)),
			4584 => std_logic_vector(to_unsigned( 158,8)),
			4585 => std_logic_vector(to_unsigned( 250,8)),
			4586 => std_logic_vector(to_unsigned( 36,8)),
			4587 => std_logic_vector(to_unsigned( 56,8)),
			4588 => std_logic_vector(to_unsigned( 219,8)),
			4589 => std_logic_vector(to_unsigned( 44,8)),
			4590 => std_logic_vector(to_unsigned( 141,8)),
			4591 => std_logic_vector(to_unsigned( 114,8)),
			4592 => std_logic_vector(to_unsigned( 85,8)),
			4593 => std_logic_vector(to_unsigned( 15,8)),
			4594 => std_logic_vector(to_unsigned( 196,8)),
			4595 => std_logic_vector(to_unsigned( 127,8)),
			4596 => std_logic_vector(to_unsigned( 248,8)),
			4597 => std_logic_vector(to_unsigned( 116,8)),
			4598 => std_logic_vector(to_unsigned( 119,8)),
			4599 => std_logic_vector(to_unsigned( 78,8)),
			4600 => std_logic_vector(to_unsigned( 171,8)),
			4601 => std_logic_vector(to_unsigned( 246,8)),
			4602 => std_logic_vector(to_unsigned( 161,8)),
			4603 => std_logic_vector(to_unsigned( 130,8)),
			4604 => std_logic_vector(to_unsigned( 169,8)),
			4605 => std_logic_vector(to_unsigned( 130,8)),
			4606 => std_logic_vector(to_unsigned( 147,8)),
			4607 => std_logic_vector(to_unsigned( 152,8)),
			4608 => std_logic_vector(to_unsigned( 156,8)),
			4609 => std_logic_vector(to_unsigned( 158,8)),
			4610 => std_logic_vector(to_unsigned( 50,8)),
			4611 => std_logic_vector(to_unsigned( 221,8)),
			4612 => std_logic_vector(to_unsigned( 53,8)),
			4613 => std_logic_vector(to_unsigned( 83,8)),
			4614 => std_logic_vector(to_unsigned( 232,8)),
			4615 => std_logic_vector(to_unsigned( 211,8)),
			4616 => std_logic_vector(to_unsigned( 93,8)),
			4617 => std_logic_vector(to_unsigned( 123,8)),
			4618 => std_logic_vector(to_unsigned( 255,8)),
			4619 => std_logic_vector(to_unsigned( 96,8)),
			4620 => std_logic_vector(to_unsigned( 211,8)),
			4621 => std_logic_vector(to_unsigned( 169,8)),
			4622 => std_logic_vector(to_unsigned( 7,8)),
			4623 => std_logic_vector(to_unsigned( 165,8)),
			4624 => std_logic_vector(to_unsigned( 210,8)),
			4625 => std_logic_vector(to_unsigned( 94,8)),
			4626 => std_logic_vector(to_unsigned( 203,8)),
			4627 => std_logic_vector(to_unsigned( 205,8)),
			4628 => std_logic_vector(to_unsigned( 214,8)),
			4629 => std_logic_vector(to_unsigned( 66,8)),
			4630 => std_logic_vector(to_unsigned( 11,8)),
			4631 => std_logic_vector(to_unsigned( 116,8)),
			4632 => std_logic_vector(to_unsigned( 158,8)),
			4633 => std_logic_vector(to_unsigned( 115,8)),
			4634 => std_logic_vector(to_unsigned( 33,8)),
			4635 => std_logic_vector(to_unsigned( 242,8)),
			4636 => std_logic_vector(to_unsigned( 125,8)),
			4637 => std_logic_vector(to_unsigned( 228,8)),
			4638 => std_logic_vector(to_unsigned( 229,8)),
			4639 => std_logic_vector(to_unsigned( 155,8)),
			4640 => std_logic_vector(to_unsigned( 91,8)),
			4641 => std_logic_vector(to_unsigned( 110,8)),
			4642 => std_logic_vector(to_unsigned( 54,8)),
			4643 => std_logic_vector(to_unsigned( 216,8)),
			4644 => std_logic_vector(to_unsigned( 92,8)),
			4645 => std_logic_vector(to_unsigned( 211,8)),
			4646 => std_logic_vector(to_unsigned( 50,8)),
			4647 => std_logic_vector(to_unsigned( 125,8)),
			4648 => std_logic_vector(to_unsigned( 194,8)),
			4649 => std_logic_vector(to_unsigned( 19,8)),
			4650 => std_logic_vector(to_unsigned( 176,8)),
			4651 => std_logic_vector(to_unsigned( 249,8)),
			4652 => std_logic_vector(to_unsigned( 254,8)),
			4653 => std_logic_vector(to_unsigned( 80,8)),
			4654 => std_logic_vector(to_unsigned( 20,8)),
			4655 => std_logic_vector(to_unsigned( 209,8)),
			4656 => std_logic_vector(to_unsigned( 149,8)),
			4657 => std_logic_vector(to_unsigned( 185,8)),
			4658 => std_logic_vector(to_unsigned( 203,8)),
			4659 => std_logic_vector(to_unsigned( 87,8)),
			4660 => std_logic_vector(to_unsigned( 241,8)),
			4661 => std_logic_vector(to_unsigned( 238,8)),
			4662 => std_logic_vector(to_unsigned( 29,8)),
			4663 => std_logic_vector(to_unsigned( 146,8)),
			4664 => std_logic_vector(to_unsigned( 74,8)),
			4665 => std_logic_vector(to_unsigned( 130,8)),
			4666 => std_logic_vector(to_unsigned( 3,8)),
			4667 => std_logic_vector(to_unsigned( 31,8)),
			4668 => std_logic_vector(to_unsigned( 37,8)),
			4669 => std_logic_vector(to_unsigned( 126,8)),
			4670 => std_logic_vector(to_unsigned( 77,8)),
			4671 => std_logic_vector(to_unsigned( 69,8)),
			4672 => std_logic_vector(to_unsigned( 189,8)),
			4673 => std_logic_vector(to_unsigned( 224,8)),
			4674 => std_logic_vector(to_unsigned( 105,8)),
			4675 => std_logic_vector(to_unsigned( 141,8)),
			4676 => std_logic_vector(to_unsigned( 123,8)),
			4677 => std_logic_vector(to_unsigned( 141,8)),
			4678 => std_logic_vector(to_unsigned( 142,8)),
			4679 => std_logic_vector(to_unsigned( 115,8)),
			4680 => std_logic_vector(to_unsigned( 183,8)),
			4681 => std_logic_vector(to_unsigned( 164,8)),
			4682 => std_logic_vector(to_unsigned( 57,8)),
			4683 => std_logic_vector(to_unsigned( 20,8)),
			4684 => std_logic_vector(to_unsigned( 221,8)),
			4685 => std_logic_vector(to_unsigned( 214,8)),
			4686 => std_logic_vector(to_unsigned( 58,8)),
			4687 => std_logic_vector(to_unsigned( 227,8)),
			4688 => std_logic_vector(to_unsigned( 172,8)),
			4689 => std_logic_vector(to_unsigned( 181,8)),
			4690 => std_logic_vector(to_unsigned( 237,8)),
			4691 => std_logic_vector(to_unsigned( 236,8)),
			4692 => std_logic_vector(to_unsigned( 200,8)),
			4693 => std_logic_vector(to_unsigned( 83,8)),
			4694 => std_logic_vector(to_unsigned( 149,8)),
			4695 => std_logic_vector(to_unsigned( 179,8)),
			4696 => std_logic_vector(to_unsigned( 84,8)),
			4697 => std_logic_vector(to_unsigned( 66,8)),
			4698 => std_logic_vector(to_unsigned( 47,8)),
			4699 => std_logic_vector(to_unsigned( 103,8)),
			4700 => std_logic_vector(to_unsigned( 230,8)),
			4701 => std_logic_vector(to_unsigned( 176,8)),
			4702 => std_logic_vector(to_unsigned( 146,8)),
			4703 => std_logic_vector(to_unsigned( 113,8)),
			4704 => std_logic_vector(to_unsigned( 191,8)),
			4705 => std_logic_vector(to_unsigned( 138,8)),
			4706 => std_logic_vector(to_unsigned( 162,8)),
			4707 => std_logic_vector(to_unsigned( 62,8)),
			4708 => std_logic_vector(to_unsigned( 174,8)),
			4709 => std_logic_vector(to_unsigned( 209,8)),
			4710 => std_logic_vector(to_unsigned( 6,8)),
			4711 => std_logic_vector(to_unsigned( 243,8)),
			4712 => std_logic_vector(to_unsigned( 129,8)),
			4713 => std_logic_vector(to_unsigned( 97,8)),
			4714 => std_logic_vector(to_unsigned( 232,8)),
			4715 => std_logic_vector(to_unsigned( 111,8)),
			4716 => std_logic_vector(to_unsigned( 185,8)),
			4717 => std_logic_vector(to_unsigned( 132,8)),
			4718 => std_logic_vector(to_unsigned( 123,8)),
			4719 => std_logic_vector(to_unsigned( 170,8)),
			4720 => std_logic_vector(to_unsigned( 230,8)),
			4721 => std_logic_vector(to_unsigned( 81,8)),
			4722 => std_logic_vector(to_unsigned( 222,8)),
			4723 => std_logic_vector(to_unsigned( 88,8)),
			4724 => std_logic_vector(to_unsigned( 233,8)),
			4725 => std_logic_vector(to_unsigned( 77,8)),
			4726 => std_logic_vector(to_unsigned( 116,8)),
			4727 => std_logic_vector(to_unsigned( 52,8)),
			4728 => std_logic_vector(to_unsigned( 229,8)),
			4729 => std_logic_vector(to_unsigned( 97,8)),
			4730 => std_logic_vector(to_unsigned( 14,8)),
			4731 => std_logic_vector(to_unsigned( 219,8)),
			4732 => std_logic_vector(to_unsigned( 229,8)),
			4733 => std_logic_vector(to_unsigned( 255,8)),
			4734 => std_logic_vector(to_unsigned( 113,8)),
			4735 => std_logic_vector(to_unsigned( 228,8)),
			4736 => std_logic_vector(to_unsigned( 123,8)),
			4737 => std_logic_vector(to_unsigned( 121,8)),
			4738 => std_logic_vector(to_unsigned( 18,8)),
			4739 => std_logic_vector(to_unsigned( 158,8)),
			4740 => std_logic_vector(to_unsigned( 252,8)),
			4741 => std_logic_vector(to_unsigned( 58,8)),
			4742 => std_logic_vector(to_unsigned( 250,8)),
			4743 => std_logic_vector(to_unsigned( 106,8)),
			4744 => std_logic_vector(to_unsigned( 119,8)),
			4745 => std_logic_vector(to_unsigned( 70,8)),
			4746 => std_logic_vector(to_unsigned( 241,8)),
			4747 => std_logic_vector(to_unsigned( 240,8)),
			4748 => std_logic_vector(to_unsigned( 84,8)),
			4749 => std_logic_vector(to_unsigned( 98,8)),
			4750 => std_logic_vector(to_unsigned( 229,8)),
			4751 => std_logic_vector(to_unsigned( 229,8)),
			4752 => std_logic_vector(to_unsigned( 19,8)),
			4753 => std_logic_vector(to_unsigned( 169,8)),
			4754 => std_logic_vector(to_unsigned( 167,8)),
			4755 => std_logic_vector(to_unsigned( 198,8)),
			4756 => std_logic_vector(to_unsigned( 24,8)),
			4757 => std_logic_vector(to_unsigned( 14,8)),
			4758 => std_logic_vector(to_unsigned( 75,8)),
			4759 => std_logic_vector(to_unsigned( 188,8)),
			4760 => std_logic_vector(to_unsigned( 101,8)),
			4761 => std_logic_vector(to_unsigned( 62,8)),
			4762 => std_logic_vector(to_unsigned( 174,8)),
			4763 => std_logic_vector(to_unsigned( 99,8)),
			4764 => std_logic_vector(to_unsigned( 102,8)),
			4765 => std_logic_vector(to_unsigned( 128,8)),
			4766 => std_logic_vector(to_unsigned( 55,8)),
			4767 => std_logic_vector(to_unsigned( 42,8)),
			4768 => std_logic_vector(to_unsigned( 98,8)),
			4769 => std_logic_vector(to_unsigned( 137,8)),
			4770 => std_logic_vector(to_unsigned( 138,8)),
			4771 => std_logic_vector(to_unsigned( 40,8)),
			4772 => std_logic_vector(to_unsigned( 34,8)),
			4773 => std_logic_vector(to_unsigned( 204,8)),
			4774 => std_logic_vector(to_unsigned( 165,8)),
			4775 => std_logic_vector(to_unsigned( 148,8)),
			4776 => std_logic_vector(to_unsigned( 235,8)),
			4777 => std_logic_vector(to_unsigned( 237,8)),
			4778 => std_logic_vector(to_unsigned( 115,8)),
			4779 => std_logic_vector(to_unsigned( 25,8)),
			4780 => std_logic_vector(to_unsigned( 171,8)),
			4781 => std_logic_vector(to_unsigned( 67,8)),
			4782 => std_logic_vector(to_unsigned( 31,8)),
			4783 => std_logic_vector(to_unsigned( 7,8)),
			4784 => std_logic_vector(to_unsigned( 4,8)),
			4785 => std_logic_vector(to_unsigned( 29,8)),
			4786 => std_logic_vector(to_unsigned( 195,8)),
			4787 => std_logic_vector(to_unsigned( 202,8)),
			4788 => std_logic_vector(to_unsigned( 220,8)),
			4789 => std_logic_vector(to_unsigned( 72,8)),
			4790 => std_logic_vector(to_unsigned( 54,8)),
			4791 => std_logic_vector(to_unsigned( 206,8)),
			4792 => std_logic_vector(to_unsigned( 233,8)),
			4793 => std_logic_vector(to_unsigned( 209,8)),
			4794 => std_logic_vector(to_unsigned( 143,8)),
			4795 => std_logic_vector(to_unsigned( 183,8)),
			4796 => std_logic_vector(to_unsigned( 143,8)),
			4797 => std_logic_vector(to_unsigned( 137,8)),
			4798 => std_logic_vector(to_unsigned( 147,8)),
			4799 => std_logic_vector(to_unsigned( 5,8)),
			4800 => std_logic_vector(to_unsigned( 77,8)),
			4801 => std_logic_vector(to_unsigned( 70,8)),
			4802 => std_logic_vector(to_unsigned( 40,8)),
			4803 => std_logic_vector(to_unsigned( 184,8)),
			4804 => std_logic_vector(to_unsigned( 99,8)),
			4805 => std_logic_vector(to_unsigned( 10,8)),
			4806 => std_logic_vector(to_unsigned( 169,8)),
			4807 => std_logic_vector(to_unsigned( 172,8)),
			4808 => std_logic_vector(to_unsigned( 47,8)),
			4809 => std_logic_vector(to_unsigned( 209,8)),
			4810 => std_logic_vector(to_unsigned( 158,8)),
			4811 => std_logic_vector(to_unsigned( 141,8)),
			4812 => std_logic_vector(to_unsigned( 61,8)),
			4813 => std_logic_vector(to_unsigned( 20,8)),
			4814 => std_logic_vector(to_unsigned( 255,8)),
			4815 => std_logic_vector(to_unsigned( 49,8)),
			4816 => std_logic_vector(to_unsigned( 154,8)),
			4817 => std_logic_vector(to_unsigned( 9,8)),
			4818 => std_logic_vector(to_unsigned( 17,8)),
			4819 => std_logic_vector(to_unsigned( 1,8)),
			4820 => std_logic_vector(to_unsigned( 1,8)),
			4821 => std_logic_vector(to_unsigned( 180,8)),
			4822 => std_logic_vector(to_unsigned( 60,8)),
			4823 => std_logic_vector(to_unsigned( 58,8)),
			4824 => std_logic_vector(to_unsigned( 162,8)),
			4825 => std_logic_vector(to_unsigned( 149,8)),
			4826 => std_logic_vector(to_unsigned( 19,8)),
			4827 => std_logic_vector(to_unsigned( 154,8)),
			4828 => std_logic_vector(to_unsigned( 160,8)),
			4829 => std_logic_vector(to_unsigned( 70,8)),
			4830 => std_logic_vector(to_unsigned( 246,8)),
			4831 => std_logic_vector(to_unsigned( 94,8)),
			4832 => std_logic_vector(to_unsigned( 229,8)),
			4833 => std_logic_vector(to_unsigned( 18,8)),
			4834 => std_logic_vector(to_unsigned( 25,8)),
			4835 => std_logic_vector(to_unsigned( 76,8)),
			4836 => std_logic_vector(to_unsigned( 219,8)),
			4837 => std_logic_vector(to_unsigned( 237,8)),
			4838 => std_logic_vector(to_unsigned( 99,8)),
			4839 => std_logic_vector(to_unsigned( 232,8)),
			4840 => std_logic_vector(to_unsigned( 32,8)),
			4841 => std_logic_vector(to_unsigned( 246,8)),
			4842 => std_logic_vector(to_unsigned( 145,8)),
			4843 => std_logic_vector(to_unsigned( 205,8)),
			4844 => std_logic_vector(to_unsigned( 218,8)),
			4845 => std_logic_vector(to_unsigned( 41,8)),
			4846 => std_logic_vector(to_unsigned( 156,8)),
			4847 => std_logic_vector(to_unsigned( 19,8)),
			4848 => std_logic_vector(to_unsigned( 107,8)),
			4849 => std_logic_vector(to_unsigned( 216,8)),
			4850 => std_logic_vector(to_unsigned( 176,8)),
			4851 => std_logic_vector(to_unsigned( 118,8)),
			4852 => std_logic_vector(to_unsigned( 108,8)),
			4853 => std_logic_vector(to_unsigned( 161,8)),
			4854 => std_logic_vector(to_unsigned( 124,8)),
			4855 => std_logic_vector(to_unsigned( 113,8)),
			4856 => std_logic_vector(to_unsigned( 88,8)),
			4857 => std_logic_vector(to_unsigned( 113,8)),
			4858 => std_logic_vector(to_unsigned( 20,8)),
			4859 => std_logic_vector(to_unsigned( 142,8)),
			4860 => std_logic_vector(to_unsigned( 203,8)),
			4861 => std_logic_vector(to_unsigned( 35,8)),
			4862 => std_logic_vector(to_unsigned( 209,8)),
			4863 => std_logic_vector(to_unsigned( 27,8)),
			4864 => std_logic_vector(to_unsigned( 143,8)),
			4865 => std_logic_vector(to_unsigned( 20,8)),
			4866 => std_logic_vector(to_unsigned( 97,8)),
			4867 => std_logic_vector(to_unsigned( 209,8)),
			4868 => std_logic_vector(to_unsigned( 70,8)),
			4869 => std_logic_vector(to_unsigned( 106,8)),
			4870 => std_logic_vector(to_unsigned( 49,8)),
			4871 => std_logic_vector(to_unsigned( 123,8)),
			4872 => std_logic_vector(to_unsigned( 108,8)),
			4873 => std_logic_vector(to_unsigned( 135,8)),
			4874 => std_logic_vector(to_unsigned( 168,8)),
			4875 => std_logic_vector(to_unsigned( 151,8)),
			4876 => std_logic_vector(to_unsigned( 19,8)),
			4877 => std_logic_vector(to_unsigned( 134,8)),
			4878 => std_logic_vector(to_unsigned( 249,8)),
			4879 => std_logic_vector(to_unsigned( 236,8)),
			4880 => std_logic_vector(to_unsigned( 4,8)),
			4881 => std_logic_vector(to_unsigned( 194,8)),
			4882 => std_logic_vector(to_unsigned( 240,8)),
			4883 => std_logic_vector(to_unsigned( 69,8)),
			4884 => std_logic_vector(to_unsigned( 6,8)),
			4885 => std_logic_vector(to_unsigned( 234,8)),
			4886 => std_logic_vector(to_unsigned( 196,8)),
			4887 => std_logic_vector(to_unsigned( 140,8)),
			4888 => std_logic_vector(to_unsigned( 31,8)),
			4889 => std_logic_vector(to_unsigned( 211,8)),
			4890 => std_logic_vector(to_unsigned( 248,8)),
			4891 => std_logic_vector(to_unsigned( 54,8)),
			4892 => std_logic_vector(to_unsigned( 162,8)),
			4893 => std_logic_vector(to_unsigned( 105,8)),
			4894 => std_logic_vector(to_unsigned( 130,8)),
			4895 => std_logic_vector(to_unsigned( 228,8)),
			4896 => std_logic_vector(to_unsigned( 83,8)),
			4897 => std_logic_vector(to_unsigned( 54,8)),
			4898 => std_logic_vector(to_unsigned( 208,8)),
			4899 => std_logic_vector(to_unsigned( 116,8)),
			4900 => std_logic_vector(to_unsigned( 184,8)),
			4901 => std_logic_vector(to_unsigned( 246,8)),
			4902 => std_logic_vector(to_unsigned( 210,8)),
			4903 => std_logic_vector(to_unsigned( 107,8)),
			4904 => std_logic_vector(to_unsigned( 78,8)),
			4905 => std_logic_vector(to_unsigned( 210,8)),
			4906 => std_logic_vector(to_unsigned( 152,8)),
			4907 => std_logic_vector(to_unsigned( 94,8)),
			4908 => std_logic_vector(to_unsigned( 120,8)),
			4909 => std_logic_vector(to_unsigned( 33,8)),
			4910 => std_logic_vector(to_unsigned( 83,8)),
			4911 => std_logic_vector(to_unsigned( 133,8)),
			4912 => std_logic_vector(to_unsigned( 224,8)),
			4913 => std_logic_vector(to_unsigned( 71,8)),
			4914 => std_logic_vector(to_unsigned( 80,8)),
			4915 => std_logic_vector(to_unsigned( 94,8)),
			4916 => std_logic_vector(to_unsigned( 90,8)),
			4917 => std_logic_vector(to_unsigned( 127,8)),
			4918 => std_logic_vector(to_unsigned( 77,8)),
			4919 => std_logic_vector(to_unsigned( 117,8)),
			4920 => std_logic_vector(to_unsigned( 66,8)),
			4921 => std_logic_vector(to_unsigned( 246,8)),
			4922 => std_logic_vector(to_unsigned( 204,8)),
			4923 => std_logic_vector(to_unsigned( 234,8)),
			4924 => std_logic_vector(to_unsigned( 78,8)),
			4925 => std_logic_vector(to_unsigned( 181,8)),
			4926 => std_logic_vector(to_unsigned( 176,8)),
			4927 => std_logic_vector(to_unsigned( 197,8)),
			4928 => std_logic_vector(to_unsigned( 224,8)),
			4929 => std_logic_vector(to_unsigned( 245,8)),
			4930 => std_logic_vector(to_unsigned( 45,8)),
			4931 => std_logic_vector(to_unsigned( 134,8)),
			4932 => std_logic_vector(to_unsigned( 88,8)),
			4933 => std_logic_vector(to_unsigned( 186,8)),
			4934 => std_logic_vector(to_unsigned( 53,8)),
			4935 => std_logic_vector(to_unsigned( 90,8)),
			4936 => std_logic_vector(to_unsigned( 92,8)),
			4937 => std_logic_vector(to_unsigned( 19,8)),
			4938 => std_logic_vector(to_unsigned( 66,8)),
			4939 => std_logic_vector(to_unsigned( 226,8)),
			4940 => std_logic_vector(to_unsigned( 45,8)),
			4941 => std_logic_vector(to_unsigned( 70,8)),
			4942 => std_logic_vector(to_unsigned( 114,8)),
			4943 => std_logic_vector(to_unsigned( 9,8)),
			4944 => std_logic_vector(to_unsigned( 198,8)),
			4945 => std_logic_vector(to_unsigned( 206,8)),
			4946 => std_logic_vector(to_unsigned( 206,8)),
			4947 => std_logic_vector(to_unsigned( 58,8)),
			4948 => std_logic_vector(to_unsigned( 231,8)),
			4949 => std_logic_vector(to_unsigned( 40,8)),
			4950 => std_logic_vector(to_unsigned( 136,8)),
			4951 => std_logic_vector(to_unsigned( 249,8)),
			4952 => std_logic_vector(to_unsigned( 242,8)),
			4953 => std_logic_vector(to_unsigned( 113,8)),
			4954 => std_logic_vector(to_unsigned( 248,8)),
			4955 => std_logic_vector(to_unsigned( 145,8)),
			4956 => std_logic_vector(to_unsigned( 85,8)),
			4957 => std_logic_vector(to_unsigned( 192,8)),
			4958 => std_logic_vector(to_unsigned( 195,8)),
			4959 => std_logic_vector(to_unsigned( 214,8)),
			4960 => std_logic_vector(to_unsigned( 242,8)),
			4961 => std_logic_vector(to_unsigned( 61,8)),
			4962 => std_logic_vector(to_unsigned( 178,8)),
			4963 => std_logic_vector(to_unsigned( 131,8)),
			4964 => std_logic_vector(to_unsigned( 83,8)),
			4965 => std_logic_vector(to_unsigned( 164,8)),
			4966 => std_logic_vector(to_unsigned( 42,8)),
			4967 => std_logic_vector(to_unsigned( 125,8)),
			4968 => std_logic_vector(to_unsigned( 18,8)),
			4969 => std_logic_vector(to_unsigned( 93,8)),
			4970 => std_logic_vector(to_unsigned( 122,8)),
			4971 => std_logic_vector(to_unsigned( 222,8)),
			4972 => std_logic_vector(to_unsigned( 245,8)),
			4973 => std_logic_vector(to_unsigned( 30,8)),
			4974 => std_logic_vector(to_unsigned( 241,8)),
			4975 => std_logic_vector(to_unsigned( 126,8)),
			4976 => std_logic_vector(to_unsigned( 186,8)),
			4977 => std_logic_vector(to_unsigned( 100,8)),
			4978 => std_logic_vector(to_unsigned( 60,8)),
			4979 => std_logic_vector(to_unsigned( 53,8)),
			4980 => std_logic_vector(to_unsigned( 21,8)),
			4981 => std_logic_vector(to_unsigned( 105,8)),
			4982 => std_logic_vector(to_unsigned( 18,8)),
			4983 => std_logic_vector(to_unsigned( 191,8)),
			4984 => std_logic_vector(to_unsigned( 56,8)),
			4985 => std_logic_vector(to_unsigned( 228,8)),
			4986 => std_logic_vector(to_unsigned( 172,8)),
			4987 => std_logic_vector(to_unsigned( 114,8)),
			4988 => std_logic_vector(to_unsigned( 99,8)),
			4989 => std_logic_vector(to_unsigned( 28,8)),
			4990 => std_logic_vector(to_unsigned( 130,8)),
			4991 => std_logic_vector(to_unsigned( 105,8)),
			4992 => std_logic_vector(to_unsigned( 13,8)),
			4993 => std_logic_vector(to_unsigned( 246,8)),
			4994 => std_logic_vector(to_unsigned( 188,8)),
			4995 => std_logic_vector(to_unsigned( 149,8)),
			4996 => std_logic_vector(to_unsigned( 210,8)),
			4997 => std_logic_vector(to_unsigned( 67,8)),
			4998 => std_logic_vector(to_unsigned( 102,8)),
			4999 => std_logic_vector(to_unsigned( 206,8)),
			5000 => std_logic_vector(to_unsigned( 23,8)),
			5001 => std_logic_vector(to_unsigned( 13,8)),
			5002 => std_logic_vector(to_unsigned( 93,8)),
			5003 => std_logic_vector(to_unsigned( 95,8)),
			5004 => std_logic_vector(to_unsigned( 45,8)),
			5005 => std_logic_vector(to_unsigned( 51,8)),
			5006 => std_logic_vector(to_unsigned( 79,8)),
			5007 => std_logic_vector(to_unsigned( 243,8)),
			5008 => std_logic_vector(to_unsigned( 22,8)),
			5009 => std_logic_vector(to_unsigned( 170,8)),
			5010 => std_logic_vector(to_unsigned( 214,8)),
			5011 => std_logic_vector(to_unsigned( 14,8)),
			5012 => std_logic_vector(to_unsigned( 63,8)),
			5013 => std_logic_vector(to_unsigned( 66,8)),
			5014 => std_logic_vector(to_unsigned( 233,8)),
			5015 => std_logic_vector(to_unsigned( 207,8)),
			5016 => std_logic_vector(to_unsigned( 167,8)),
			5017 => std_logic_vector(to_unsigned( 63,8)),
			5018 => std_logic_vector(to_unsigned( 126,8)),
			5019 => std_logic_vector(to_unsigned( 219,8)),
			5020 => std_logic_vector(to_unsigned( 131,8)),
			5021 => std_logic_vector(to_unsigned( 205,8)),
			5022 => std_logic_vector(to_unsigned( 44,8)),
			5023 => std_logic_vector(to_unsigned( 116,8)),
			5024 => std_logic_vector(to_unsigned( 96,8)),
			5025 => std_logic_vector(to_unsigned( 224,8)),
			5026 => std_logic_vector(to_unsigned( 40,8)),
			5027 => std_logic_vector(to_unsigned( 37,8)),
			5028 => std_logic_vector(to_unsigned( 192,8)),
			5029 => std_logic_vector(to_unsigned( 21,8)),
			5030 => std_logic_vector(to_unsigned( 166,8)),
			5031 => std_logic_vector(to_unsigned( 151,8)),
			5032 => std_logic_vector(to_unsigned( 10,8)),
			5033 => std_logic_vector(to_unsigned( 172,8)),
			5034 => std_logic_vector(to_unsigned( 90,8)),
			5035 => std_logic_vector(to_unsigned( 109,8)),
			5036 => std_logic_vector(to_unsigned( 45,8)),
			5037 => std_logic_vector(to_unsigned( 119,8)),
			5038 => std_logic_vector(to_unsigned( 0,8)),
			5039 => std_logic_vector(to_unsigned( 81,8)),
			5040 => std_logic_vector(to_unsigned( 214,8)),
			5041 => std_logic_vector(to_unsigned( 96,8)),
			5042 => std_logic_vector(to_unsigned( 95,8)),
			5043 => std_logic_vector(to_unsigned( 59,8)),
			5044 => std_logic_vector(to_unsigned( 239,8)),
			5045 => std_logic_vector(to_unsigned( 155,8)),
			5046 => std_logic_vector(to_unsigned( 217,8)),
			5047 => std_logic_vector(to_unsigned( 161,8)),
			5048 => std_logic_vector(to_unsigned( 46,8)),
			5049 => std_logic_vector(to_unsigned( 29,8)),
			5050 => std_logic_vector(to_unsigned( 236,8)),
			5051 => std_logic_vector(to_unsigned( 163,8)),
			5052 => std_logic_vector(to_unsigned( 137,8)),
			5053 => std_logic_vector(to_unsigned( 31,8)),
			5054 => std_logic_vector(to_unsigned( 55,8)),
			5055 => std_logic_vector(to_unsigned( 24,8)),
			5056 => std_logic_vector(to_unsigned( 236,8)),
			5057 => std_logic_vector(to_unsigned( 144,8)),
			5058 => std_logic_vector(to_unsigned( 199,8)),
			5059 => std_logic_vector(to_unsigned( 158,8)),
			5060 => std_logic_vector(to_unsigned( 35,8)),
			5061 => std_logic_vector(to_unsigned( 141,8)),
			5062 => std_logic_vector(to_unsigned( 173,8)),
			5063 => std_logic_vector(to_unsigned( 154,8)),
			5064 => std_logic_vector(to_unsigned( 5,8)),
			5065 => std_logic_vector(to_unsigned( 19,8)),
			5066 => std_logic_vector(to_unsigned( 253,8)),
			5067 => std_logic_vector(to_unsigned( 46,8)),
			5068 => std_logic_vector(to_unsigned( 68,8)),
			5069 => std_logic_vector(to_unsigned( 168,8)),
			5070 => std_logic_vector(to_unsigned( 21,8)),
			5071 => std_logic_vector(to_unsigned( 101,8)),
			5072 => std_logic_vector(to_unsigned( 188,8)),
			5073 => std_logic_vector(to_unsigned( 107,8)),
			5074 => std_logic_vector(to_unsigned( 17,8)),
			5075 => std_logic_vector(to_unsigned( 165,8)),
			5076 => std_logic_vector(to_unsigned( 227,8)),
			5077 => std_logic_vector(to_unsigned( 253,8)),
			5078 => std_logic_vector(to_unsigned( 8,8)),
			5079 => std_logic_vector(to_unsigned( 91,8)),
			5080 => std_logic_vector(to_unsigned( 171,8)),
			5081 => std_logic_vector(to_unsigned( 31,8)),
			5082 => std_logic_vector(to_unsigned( 4,8)),
			5083 => std_logic_vector(to_unsigned( 112,8)),
			5084 => std_logic_vector(to_unsigned( 156,8)),
			5085 => std_logic_vector(to_unsigned( 151,8)),
			5086 => std_logic_vector(to_unsigned( 247,8)),
			5087 => std_logic_vector(to_unsigned( 231,8)),
			5088 => std_logic_vector(to_unsigned( 143,8)),
			5089 => std_logic_vector(to_unsigned( 174,8)),
			5090 => std_logic_vector(to_unsigned( 150,8)),
			5091 => std_logic_vector(to_unsigned( 77,8)),
			5092 => std_logic_vector(to_unsigned( 14,8)),
			5093 => std_logic_vector(to_unsigned( 172,8)),
			5094 => std_logic_vector(to_unsigned( 129,8)),
			5095 => std_logic_vector(to_unsigned( 125,8)),
			5096 => std_logic_vector(to_unsigned( 208,8)),
			5097 => std_logic_vector(to_unsigned( 249,8)),
			5098 => std_logic_vector(to_unsigned( 138,8)),
			5099 => std_logic_vector(to_unsigned( 100,8)),
			5100 => std_logic_vector(to_unsigned( 183,8)),
			5101 => std_logic_vector(to_unsigned( 248,8)),
			5102 => std_logic_vector(to_unsigned( 82,8)),
			5103 => std_logic_vector(to_unsigned( 59,8)),
			5104 => std_logic_vector(to_unsigned( 137,8)),
			5105 => std_logic_vector(to_unsigned( 190,8)),
			5106 => std_logic_vector(to_unsigned( 18,8)),
			5107 => std_logic_vector(to_unsigned( 153,8)),
			5108 => std_logic_vector(to_unsigned( 251,8)),
			5109 => std_logic_vector(to_unsigned( 236,8)),
			5110 => std_logic_vector(to_unsigned( 104,8)),
			5111 => std_logic_vector(to_unsigned( 46,8)),
			5112 => std_logic_vector(to_unsigned( 239,8)),
			5113 => std_logic_vector(to_unsigned( 200,8)),
			5114 => std_logic_vector(to_unsigned( 128,8)),
			5115 => std_logic_vector(to_unsigned( 158,8)),
			5116 => std_logic_vector(to_unsigned( 106,8)),
			5117 => std_logic_vector(to_unsigned( 202,8)),
			5118 => std_logic_vector(to_unsigned( 91,8)),
			5119 => std_logic_vector(to_unsigned( 174,8)),
			5120 => std_logic_vector(to_unsigned( 87,8)),
			5121 => std_logic_vector(to_unsigned( 192,8)),
			5122 => std_logic_vector(to_unsigned( 215,8)),
			5123 => std_logic_vector(to_unsigned( 16,8)),
			5124 => std_logic_vector(to_unsigned( 200,8)),
			5125 => std_logic_vector(to_unsigned( 161,8)),
			5126 => std_logic_vector(to_unsigned( 103,8)),
			5127 => std_logic_vector(to_unsigned( 75,8)),
			5128 => std_logic_vector(to_unsigned( 121,8)),
			5129 => std_logic_vector(to_unsigned( 24,8)),
			5130 => std_logic_vector(to_unsigned( 5,8)),
			5131 => std_logic_vector(to_unsigned( 56,8)),
			5132 => std_logic_vector(to_unsigned( 153,8)),
			5133 => std_logic_vector(to_unsigned( 142,8)),
			5134 => std_logic_vector(to_unsigned( 17,8)),
			5135 => std_logic_vector(to_unsigned( 79,8)),
			5136 => std_logic_vector(to_unsigned( 148,8)),
			5137 => std_logic_vector(to_unsigned( 29,8)),
			5138 => std_logic_vector(to_unsigned( 59,8)),
			5139 => std_logic_vector(to_unsigned( 57,8)),
			5140 => std_logic_vector(to_unsigned( 32,8)),
			5141 => std_logic_vector(to_unsigned( 41,8)),
			5142 => std_logic_vector(to_unsigned( 150,8)),
			5143 => std_logic_vector(to_unsigned( 157,8)),
			5144 => std_logic_vector(to_unsigned( 35,8)),
			5145 => std_logic_vector(to_unsigned( 185,8)),
			5146 => std_logic_vector(to_unsigned( 195,8)),
			5147 => std_logic_vector(to_unsigned( 2,8)),
			5148 => std_logic_vector(to_unsigned( 103,8)),
			5149 => std_logic_vector(to_unsigned( 92,8)),
			5150 => std_logic_vector(to_unsigned( 164,8)),
			5151 => std_logic_vector(to_unsigned( 11,8)),
			5152 => std_logic_vector(to_unsigned( 219,8)),
			5153 => std_logic_vector(to_unsigned( 214,8)),
			5154 => std_logic_vector(to_unsigned( 238,8)),
			5155 => std_logic_vector(to_unsigned( 107,8)),
			5156 => std_logic_vector(to_unsigned( 38,8)),
			5157 => std_logic_vector(to_unsigned( 29,8)),
			5158 => std_logic_vector(to_unsigned( 250,8)),
			5159 => std_logic_vector(to_unsigned( 58,8)),
			5160 => std_logic_vector(to_unsigned( 87,8)),
			5161 => std_logic_vector(to_unsigned( 70,8)),
			5162 => std_logic_vector(to_unsigned( 163,8)),
			5163 => std_logic_vector(to_unsigned( 183,8)),
			5164 => std_logic_vector(to_unsigned( 77,8)),
			5165 => std_logic_vector(to_unsigned( 235,8)),
			5166 => std_logic_vector(to_unsigned( 72,8)),
			5167 => std_logic_vector(to_unsigned( 227,8)),
			5168 => std_logic_vector(to_unsigned( 59,8)),
			5169 => std_logic_vector(to_unsigned( 40,8)),
			5170 => std_logic_vector(to_unsigned( 86,8)),
			5171 => std_logic_vector(to_unsigned( 144,8)),
			5172 => std_logic_vector(to_unsigned( 178,8)),
			5173 => std_logic_vector(to_unsigned( 59,8)),
			5174 => std_logic_vector(to_unsigned( 254,8)),
			5175 => std_logic_vector(to_unsigned( 190,8)),
			5176 => std_logic_vector(to_unsigned( 85,8)),
			5177 => std_logic_vector(to_unsigned( 3,8)),
			5178 => std_logic_vector(to_unsigned( 145,8)),
			5179 => std_logic_vector(to_unsigned( 196,8)),
			5180 => std_logic_vector(to_unsigned( 60,8)),
			5181 => std_logic_vector(to_unsigned( 26,8)),
			5182 => std_logic_vector(to_unsigned( 255,8)),
			5183 => std_logic_vector(to_unsigned( 49,8)),
			5184 => std_logic_vector(to_unsigned( 219,8)),
			5185 => std_logic_vector(to_unsigned( 8,8)),
			5186 => std_logic_vector(to_unsigned( 77,8)),
			5187 => std_logic_vector(to_unsigned( 253,8)),
			5188 => std_logic_vector(to_unsigned( 0,8)),
			5189 => std_logic_vector(to_unsigned( 253,8)),
			5190 => std_logic_vector(to_unsigned( 223,8)),
			5191 => std_logic_vector(to_unsigned( 106,8)),
			5192 => std_logic_vector(to_unsigned( 14,8)),
			5193 => std_logic_vector(to_unsigned( 206,8)),
			5194 => std_logic_vector(to_unsigned( 125,8)),
			5195 => std_logic_vector(to_unsigned( 211,8)),
			5196 => std_logic_vector(to_unsigned( 235,8)),
			5197 => std_logic_vector(to_unsigned( 15,8)),
			5198 => std_logic_vector(to_unsigned( 236,8)),
			5199 => std_logic_vector(to_unsigned( 134,8)),
			5200 => std_logic_vector(to_unsigned( 43,8)),
			5201 => std_logic_vector(to_unsigned( 147,8)),
			5202 => std_logic_vector(to_unsigned( 139,8)),
			5203 => std_logic_vector(to_unsigned( 67,8)),
			5204 => std_logic_vector(to_unsigned( 48,8)),
			5205 => std_logic_vector(to_unsigned( 26,8)),
			5206 => std_logic_vector(to_unsigned( 212,8)),
			5207 => std_logic_vector(to_unsigned( 158,8)),
			5208 => std_logic_vector(to_unsigned( 21,8)),
			5209 => std_logic_vector(to_unsigned( 199,8)),
			5210 => std_logic_vector(to_unsigned( 233,8)),
			5211 => std_logic_vector(to_unsigned( 213,8)),
			5212 => std_logic_vector(to_unsigned( 228,8)),
			5213 => std_logic_vector(to_unsigned( 234,8)),
			5214 => std_logic_vector(to_unsigned( 3,8)),
			5215 => std_logic_vector(to_unsigned( 7,8)),
			5216 => std_logic_vector(to_unsigned( 210,8)),
			5217 => std_logic_vector(to_unsigned( 97,8)),
			5218 => std_logic_vector(to_unsigned( 50,8)),
			5219 => std_logic_vector(to_unsigned( 184,8)),
			5220 => std_logic_vector(to_unsigned( 188,8)),
			5221 => std_logic_vector(to_unsigned( 240,8)),
			5222 => std_logic_vector(to_unsigned( 144,8)),
			5223 => std_logic_vector(to_unsigned( 97,8)),
			5224 => std_logic_vector(to_unsigned( 41,8)),
			5225 => std_logic_vector(to_unsigned( 99,8)),
			5226 => std_logic_vector(to_unsigned( 14,8)),
			5227 => std_logic_vector(to_unsigned( 155,8)),
			5228 => std_logic_vector(to_unsigned( 5,8)),
			5229 => std_logic_vector(to_unsigned( 111,8)),
			5230 => std_logic_vector(to_unsigned( 216,8)),
			5231 => std_logic_vector(to_unsigned( 156,8)),
			5232 => std_logic_vector(to_unsigned( 158,8)),
			5233 => std_logic_vector(to_unsigned( 137,8)),
			5234 => std_logic_vector(to_unsigned( 88,8)),
			5235 => std_logic_vector(to_unsigned( 107,8)),
			5236 => std_logic_vector(to_unsigned( 105,8)),
			5237 => std_logic_vector(to_unsigned( 162,8)),
			5238 => std_logic_vector(to_unsigned( 187,8)),
			5239 => std_logic_vector(to_unsigned( 248,8)),
			5240 => std_logic_vector(to_unsigned( 67,8)),
			5241 => std_logic_vector(to_unsigned( 185,8)),
			5242 => std_logic_vector(to_unsigned( 5,8)),
			5243 => std_logic_vector(to_unsigned( 15,8)),
			5244 => std_logic_vector(to_unsigned( 158,8)),
			5245 => std_logic_vector(to_unsigned( 111,8)),
			5246 => std_logic_vector(to_unsigned( 149,8)),
			5247 => std_logic_vector(to_unsigned( 40,8)),
			5248 => std_logic_vector(to_unsigned( 25,8)),
			5249 => std_logic_vector(to_unsigned( 145,8)),
			5250 => std_logic_vector(to_unsigned( 209,8)),
			5251 => std_logic_vector(to_unsigned( 246,8)),
			5252 => std_logic_vector(to_unsigned( 9,8)),
			5253 => std_logic_vector(to_unsigned( 180,8)),
			5254 => std_logic_vector(to_unsigned( 176,8)),
			5255 => std_logic_vector(to_unsigned( 44,8)),
			5256 => std_logic_vector(to_unsigned( 217,8)),
			5257 => std_logic_vector(to_unsigned( 201,8)),
			5258 => std_logic_vector(to_unsigned( 171,8)),
			5259 => std_logic_vector(to_unsigned( 141,8)),
			5260 => std_logic_vector(to_unsigned( 34,8)),
			5261 => std_logic_vector(to_unsigned( 50,8)),
			5262 => std_logic_vector(to_unsigned( 178,8)),
			5263 => std_logic_vector(to_unsigned( 113,8)),
			5264 => std_logic_vector(to_unsigned( 196,8)),
			5265 => std_logic_vector(to_unsigned( 171,8)),
			5266 => std_logic_vector(to_unsigned( 124,8)),
			5267 => std_logic_vector(to_unsigned( 108,8)),
			5268 => std_logic_vector(to_unsigned( 228,8)),
			5269 => std_logic_vector(to_unsigned( 190,8)),
			5270 => std_logic_vector(to_unsigned( 110,8)),
			5271 => std_logic_vector(to_unsigned( 88,8)),
			5272 => std_logic_vector(to_unsigned( 82,8)),
			5273 => std_logic_vector(to_unsigned( 19,8)),
			5274 => std_logic_vector(to_unsigned( 24,8)),
			5275 => std_logic_vector(to_unsigned( 10,8)),
			5276 => std_logic_vector(to_unsigned( 167,8)),
			5277 => std_logic_vector(to_unsigned( 59,8)),
			5278 => std_logic_vector(to_unsigned( 181,8)),
			5279 => std_logic_vector(to_unsigned( 133,8)),
			5280 => std_logic_vector(to_unsigned( 63,8)),
			5281 => std_logic_vector(to_unsigned( 103,8)),
			5282 => std_logic_vector(to_unsigned( 5,8)),
			5283 => std_logic_vector(to_unsigned( 239,8)),
			5284 => std_logic_vector(to_unsigned( 222,8)),
			5285 => std_logic_vector(to_unsigned( 12,8)),
			5286 => std_logic_vector(to_unsigned( 130,8)),
			5287 => std_logic_vector(to_unsigned( 246,8)),
			5288 => std_logic_vector(to_unsigned( 3,8)),
			5289 => std_logic_vector(to_unsigned( 108,8)),
			5290 => std_logic_vector(to_unsigned( 97,8)),
			5291 => std_logic_vector(to_unsigned( 250,8)),
			5292 => std_logic_vector(to_unsigned( 117,8)),
			5293 => std_logic_vector(to_unsigned( 175,8)),
			5294 => std_logic_vector(to_unsigned( 219,8)),
			5295 => std_logic_vector(to_unsigned( 192,8)),
			5296 => std_logic_vector(to_unsigned( 178,8)),
			5297 => std_logic_vector(to_unsigned( 10,8)),
			5298 => std_logic_vector(to_unsigned( 114,8)),
			5299 => std_logic_vector(to_unsigned( 45,8)),
			5300 => std_logic_vector(to_unsigned( 107,8)),
			5301 => std_logic_vector(to_unsigned( 109,8)),
			5302 => std_logic_vector(to_unsigned( 1,8)),
			5303 => std_logic_vector(to_unsigned( 104,8)),
			5304 => std_logic_vector(to_unsigned( 96,8)),
			5305 => std_logic_vector(to_unsigned( 157,8)),
			5306 => std_logic_vector(to_unsigned( 209,8)),
			5307 => std_logic_vector(to_unsigned( 122,8)),
			5308 => std_logic_vector(to_unsigned( 20,8)),
			5309 => std_logic_vector(to_unsigned( 34,8)),
			5310 => std_logic_vector(to_unsigned( 156,8)),
			5311 => std_logic_vector(to_unsigned( 238,8)),
			5312 => std_logic_vector(to_unsigned( 114,8)),
			5313 => std_logic_vector(to_unsigned( 241,8)),
			5314 => std_logic_vector(to_unsigned( 246,8)),
			5315 => std_logic_vector(to_unsigned( 159,8)),
			5316 => std_logic_vector(to_unsigned( 147,8)),
			5317 => std_logic_vector(to_unsigned( 161,8)),
			5318 => std_logic_vector(to_unsigned( 80,8)),
			5319 => std_logic_vector(to_unsigned( 72,8)),
			5320 => std_logic_vector(to_unsigned( 82,8)),
			5321 => std_logic_vector(to_unsigned( 83,8)),
			5322 => std_logic_vector(to_unsigned( 27,8)),
			5323 => std_logic_vector(to_unsigned( 244,8)),
			5324 => std_logic_vector(to_unsigned( 203,8)),
			5325 => std_logic_vector(to_unsigned( 253,8)),
			5326 => std_logic_vector(to_unsigned( 0,8)),
			5327 => std_logic_vector(to_unsigned( 30,8)),
			5328 => std_logic_vector(to_unsigned( 207,8)),
			5329 => std_logic_vector(to_unsigned( 191,8)),
			5330 => std_logic_vector(to_unsigned( 142,8)),
			5331 => std_logic_vector(to_unsigned( 13,8)),
			5332 => std_logic_vector(to_unsigned( 172,8)),
			5333 => std_logic_vector(to_unsigned( 135,8)),
			5334 => std_logic_vector(to_unsigned( 107,8)),
			5335 => std_logic_vector(to_unsigned( 182,8)),
			5336 => std_logic_vector(to_unsigned( 11,8)),
			5337 => std_logic_vector(to_unsigned( 87,8)),
			5338 => std_logic_vector(to_unsigned( 143,8)),
			5339 => std_logic_vector(to_unsigned( 115,8)),
			5340 => std_logic_vector(to_unsigned( 230,8)),
			5341 => std_logic_vector(to_unsigned( 210,8)),
			5342 => std_logic_vector(to_unsigned( 64,8)),
			5343 => std_logic_vector(to_unsigned( 40,8)),
			5344 => std_logic_vector(to_unsigned( 119,8)),
			5345 => std_logic_vector(to_unsigned( 114,8)),
			5346 => std_logic_vector(to_unsigned( 68,8)),
			5347 => std_logic_vector(to_unsigned( 208,8)),
			5348 => std_logic_vector(to_unsigned( 81,8)),
			5349 => std_logic_vector(to_unsigned( 219,8)),
			5350 => std_logic_vector(to_unsigned( 36,8)),
			5351 => std_logic_vector(to_unsigned( 73,8)),
			5352 => std_logic_vector(to_unsigned( 139,8)),
			5353 => std_logic_vector(to_unsigned( 125,8)),
			5354 => std_logic_vector(to_unsigned( 77,8)),
			5355 => std_logic_vector(to_unsigned( 100,8)),
			5356 => std_logic_vector(to_unsigned( 161,8)),
			5357 => std_logic_vector(to_unsigned( 10,8)),
			5358 => std_logic_vector(to_unsigned( 197,8)),
			5359 => std_logic_vector(to_unsigned( 169,8)),
			5360 => std_logic_vector(to_unsigned( 63,8)),
			5361 => std_logic_vector(to_unsigned( 222,8)),
			5362 => std_logic_vector(to_unsigned( 153,8)),
			5363 => std_logic_vector(to_unsigned( 223,8)),
			5364 => std_logic_vector(to_unsigned( 45,8)),
			5365 => std_logic_vector(to_unsigned( 73,8)),
			5366 => std_logic_vector(to_unsigned( 243,8)),
			5367 => std_logic_vector(to_unsigned( 222,8)),
			5368 => std_logic_vector(to_unsigned( 214,8)),
			5369 => std_logic_vector(to_unsigned( 3,8)),
			5370 => std_logic_vector(to_unsigned( 140,8)),
			5371 => std_logic_vector(to_unsigned( 209,8)),
			5372 => std_logic_vector(to_unsigned( 145,8)),
			5373 => std_logic_vector(to_unsigned( 251,8)),
			5374 => std_logic_vector(to_unsigned( 0,8)),
			5375 => std_logic_vector(to_unsigned( 50,8)),
			5376 => std_logic_vector(to_unsigned( 43,8)),
			5377 => std_logic_vector(to_unsigned( 88,8)),
			5378 => std_logic_vector(to_unsigned( 200,8)),
			5379 => std_logic_vector(to_unsigned( 146,8)),
			5380 => std_logic_vector(to_unsigned( 192,8)),
			5381 => std_logic_vector(to_unsigned( 184,8)),
			5382 => std_logic_vector(to_unsigned( 33,8)),
			5383 => std_logic_vector(to_unsigned( 198,8)),
			5384 => std_logic_vector(to_unsigned( 180,8)),
			5385 => std_logic_vector(to_unsigned( 178,8)),
			5386 => std_logic_vector(to_unsigned( 4,8)),
			5387 => std_logic_vector(to_unsigned( 166,8)),
			5388 => std_logic_vector(to_unsigned( 209,8)),
			5389 => std_logic_vector(to_unsigned( 192,8)),
			5390 => std_logic_vector(to_unsigned( 158,8)),
			5391 => std_logic_vector(to_unsigned( 246,8)),
			5392 => std_logic_vector(to_unsigned( 111,8)),
			5393 => std_logic_vector(to_unsigned( 32,8)),
			5394 => std_logic_vector(to_unsigned( 31,8)),
			5395 => std_logic_vector(to_unsigned( 215,8)),
			5396 => std_logic_vector(to_unsigned( 246,8)),
			5397 => std_logic_vector(to_unsigned( 249,8)),
			5398 => std_logic_vector(to_unsigned( 28,8)),
			5399 => std_logic_vector(to_unsigned( 55,8)),
			5400 => std_logic_vector(to_unsigned( 145,8)),
			5401 => std_logic_vector(to_unsigned( 190,8)),
			5402 => std_logic_vector(to_unsigned( 130,8)),
			5403 => std_logic_vector(to_unsigned( 246,8)),
			5404 => std_logic_vector(to_unsigned( 9,8)),
			5405 => std_logic_vector(to_unsigned( 160,8)),
			5406 => std_logic_vector(to_unsigned( 25,8)),
			5407 => std_logic_vector(to_unsigned( 153,8)),
			5408 => std_logic_vector(to_unsigned( 181,8)),
			5409 => std_logic_vector(to_unsigned( 214,8)),
			5410 => std_logic_vector(to_unsigned( 80,8)),
			5411 => std_logic_vector(to_unsigned( 184,8)),
			5412 => std_logic_vector(to_unsigned( 138,8)),
			5413 => std_logic_vector(to_unsigned( 2,8)),
			5414 => std_logic_vector(to_unsigned( 44,8)),
			5415 => std_logic_vector(to_unsigned( 9,8)),
			5416 => std_logic_vector(to_unsigned( 240,8)),
			5417 => std_logic_vector(to_unsigned( 176,8)),
			5418 => std_logic_vector(to_unsigned( 60,8)),
			5419 => std_logic_vector(to_unsigned( 117,8)),
			5420 => std_logic_vector(to_unsigned( 195,8)),
			5421 => std_logic_vector(to_unsigned( 135,8)),
			5422 => std_logic_vector(to_unsigned( 227,8)),
			5423 => std_logic_vector(to_unsigned( 230,8)),
			5424 => std_logic_vector(to_unsigned( 82,8)),
			5425 => std_logic_vector(to_unsigned( 79,8)),
			5426 => std_logic_vector(to_unsigned( 241,8)),
			5427 => std_logic_vector(to_unsigned( 243,8)),
			5428 => std_logic_vector(to_unsigned( 44,8)),
			5429 => std_logic_vector(to_unsigned( 113,8)),
			5430 => std_logic_vector(to_unsigned( 81,8)),
			5431 => std_logic_vector(to_unsigned( 25,8)),
			5432 => std_logic_vector(to_unsigned( 118,8)),
			5433 => std_logic_vector(to_unsigned( 191,8)),
			5434 => std_logic_vector(to_unsigned( 165,8)),
			5435 => std_logic_vector(to_unsigned( 37,8)),
			5436 => std_logic_vector(to_unsigned( 87,8)),
			5437 => std_logic_vector(to_unsigned( 208,8)),
			5438 => std_logic_vector(to_unsigned( 252,8)),
			5439 => std_logic_vector(to_unsigned( 233,8)),
			5440 => std_logic_vector(to_unsigned( 251,8)),
			5441 => std_logic_vector(to_unsigned( 219,8)),
			5442 => std_logic_vector(to_unsigned( 103,8)),
			5443 => std_logic_vector(to_unsigned( 248,8)),
			5444 => std_logic_vector(to_unsigned( 242,8)),
			5445 => std_logic_vector(to_unsigned( 113,8)),
			5446 => std_logic_vector(to_unsigned( 128,8)),
			5447 => std_logic_vector(to_unsigned( 91,8)),
			5448 => std_logic_vector(to_unsigned( 214,8)),
			5449 => std_logic_vector(to_unsigned( 209,8)),
			5450 => std_logic_vector(to_unsigned( 95,8)),
			5451 => std_logic_vector(to_unsigned( 138,8)),
			5452 => std_logic_vector(to_unsigned( 180,8)),
			5453 => std_logic_vector(to_unsigned( 164,8)),
			5454 => std_logic_vector(to_unsigned( 243,8)),
			5455 => std_logic_vector(to_unsigned( 121,8)),
			5456 => std_logic_vector(to_unsigned( 126,8)),
			5457 => std_logic_vector(to_unsigned( 98,8)),
			5458 => std_logic_vector(to_unsigned( 44,8)),
			5459 => std_logic_vector(to_unsigned( 187,8)),
			5460 => std_logic_vector(to_unsigned( 61,8)),
			5461 => std_logic_vector(to_unsigned( 172,8)),
			5462 => std_logic_vector(to_unsigned( 168,8)),
			5463 => std_logic_vector(to_unsigned( 37,8)),
			5464 => std_logic_vector(to_unsigned( 68,8)),
			5465 => std_logic_vector(to_unsigned( 12,8)),
			5466 => std_logic_vector(to_unsigned( 248,8)),
			5467 => std_logic_vector(to_unsigned( 3,8)),
			5468 => std_logic_vector(to_unsigned( 183,8)),
			5469 => std_logic_vector(to_unsigned( 132,8)),
			5470 => std_logic_vector(to_unsigned( 226,8)),
			5471 => std_logic_vector(to_unsigned( 21,8)),
			5472 => std_logic_vector(to_unsigned( 167,8)),
			5473 => std_logic_vector(to_unsigned( 205,8)),
			5474 => std_logic_vector(to_unsigned( 162,8)),
			5475 => std_logic_vector(to_unsigned( 237,8)),
			5476 => std_logic_vector(to_unsigned( 22,8)),
			5477 => std_logic_vector(to_unsigned( 113,8)),
			5478 => std_logic_vector(to_unsigned( 96,8)),
			5479 => std_logic_vector(to_unsigned( 78,8)),
			5480 => std_logic_vector(to_unsigned( 192,8)),
			5481 => std_logic_vector(to_unsigned( 102,8)),
			5482 => std_logic_vector(to_unsigned( 141,8)),
			5483 => std_logic_vector(to_unsigned( 222,8)),
			5484 => std_logic_vector(to_unsigned( 127,8)),
			5485 => std_logic_vector(to_unsigned( 14,8)),
			5486 => std_logic_vector(to_unsigned( 210,8)),
			5487 => std_logic_vector(to_unsigned( 86,8)),
			5488 => std_logic_vector(to_unsigned( 148,8)),
			5489 => std_logic_vector(to_unsigned( 174,8)),
			5490 => std_logic_vector(to_unsigned( 37,8)),
			5491 => std_logic_vector(to_unsigned( 157,8)),
			5492 => std_logic_vector(to_unsigned( 75,8)),
			5493 => std_logic_vector(to_unsigned( 127,8)),
			5494 => std_logic_vector(to_unsigned( 239,8)),
			5495 => std_logic_vector(to_unsigned( 102,8)),
			5496 => std_logic_vector(to_unsigned( 45,8)),
			5497 => std_logic_vector(to_unsigned( 96,8)),
			5498 => std_logic_vector(to_unsigned( 117,8)),
			5499 => std_logic_vector(to_unsigned( 79,8)),
			5500 => std_logic_vector(to_unsigned( 113,8)),
			5501 => std_logic_vector(to_unsigned( 189,8)),
			5502 => std_logic_vector(to_unsigned( 41,8)),
			5503 => std_logic_vector(to_unsigned( 134,8)),
			5504 => std_logic_vector(to_unsigned( 132,8)),
			5505 => std_logic_vector(to_unsigned( 35,8)),
			5506 => std_logic_vector(to_unsigned( 91,8)),
			5507 => std_logic_vector(to_unsigned( 157,8)),
			5508 => std_logic_vector(to_unsigned( 86,8)),
			5509 => std_logic_vector(to_unsigned( 219,8)),
			5510 => std_logic_vector(to_unsigned( 50,8)),
			5511 => std_logic_vector(to_unsigned( 84,8)),
			5512 => std_logic_vector(to_unsigned( 153,8)),
			5513 => std_logic_vector(to_unsigned( 13,8)),
			5514 => std_logic_vector(to_unsigned( 63,8)),
			5515 => std_logic_vector(to_unsigned( 33,8)),
			5516 => std_logic_vector(to_unsigned( 15,8)),
			5517 => std_logic_vector(to_unsigned( 228,8)),
			5518 => std_logic_vector(to_unsigned( 28,8)),
			5519 => std_logic_vector(to_unsigned( 184,8)),
			5520 => std_logic_vector(to_unsigned( 33,8)),
			5521 => std_logic_vector(to_unsigned( 38,8)),
			5522 => std_logic_vector(to_unsigned( 208,8)),
			5523 => std_logic_vector(to_unsigned( 187,8)),
			5524 => std_logic_vector(to_unsigned( 33,8)),
			5525 => std_logic_vector(to_unsigned( 24,8)),
			5526 => std_logic_vector(to_unsigned( 148,8)),
			5527 => std_logic_vector(to_unsigned( 199,8)),
			5528 => std_logic_vector(to_unsigned( 191,8)),
			5529 => std_logic_vector(to_unsigned( 35,8)),
			5530 => std_logic_vector(to_unsigned( 95,8)),
			5531 => std_logic_vector(to_unsigned( 215,8)),
			5532 => std_logic_vector(to_unsigned( 191,8)),
			5533 => std_logic_vector(to_unsigned( 245,8)),
			5534 => std_logic_vector(to_unsigned( 106,8)),
			5535 => std_logic_vector(to_unsigned( 135,8)),
			5536 => std_logic_vector(to_unsigned( 41,8)),
			5537 => std_logic_vector(to_unsigned( 115,8)),
			5538 => std_logic_vector(to_unsigned( 140,8)),
			5539 => std_logic_vector(to_unsigned( 130,8)),
			5540 => std_logic_vector(to_unsigned( 11,8)),
			5541 => std_logic_vector(to_unsigned( 66,8)),
			5542 => std_logic_vector(to_unsigned( 236,8)),
			5543 => std_logic_vector(to_unsigned( 125,8)),
			5544 => std_logic_vector(to_unsigned( 63,8)),
			5545 => std_logic_vector(to_unsigned( 116,8)),
			5546 => std_logic_vector(to_unsigned( 195,8)),
			5547 => std_logic_vector(to_unsigned( 247,8)),
			5548 => std_logic_vector(to_unsigned( 96,8)),
			5549 => std_logic_vector(to_unsigned( 169,8)),
			5550 => std_logic_vector(to_unsigned( 146,8)),
			5551 => std_logic_vector(to_unsigned( 220,8)),
			5552 => std_logic_vector(to_unsigned( 124,8)),
			5553 => std_logic_vector(to_unsigned( 88,8)),
			5554 => std_logic_vector(to_unsigned( 41,8)),
			5555 => std_logic_vector(to_unsigned( 182,8)),
			5556 => std_logic_vector(to_unsigned( 176,8)),
			5557 => std_logic_vector(to_unsigned( 113,8)),
			5558 => std_logic_vector(to_unsigned( 68,8)),
			5559 => std_logic_vector(to_unsigned( 9,8)),
			5560 => std_logic_vector(to_unsigned( 250,8)),
			5561 => std_logic_vector(to_unsigned( 79,8)),
			5562 => std_logic_vector(to_unsigned( 53,8)),
			5563 => std_logic_vector(to_unsigned( 247,8)),
			5564 => std_logic_vector(to_unsigned( 216,8)),
			5565 => std_logic_vector(to_unsigned( 76,8)),
			5566 => std_logic_vector(to_unsigned( 142,8)),
			5567 => std_logic_vector(to_unsigned( 176,8)),
			5568 => std_logic_vector(to_unsigned( 100,8)),
			5569 => std_logic_vector(to_unsigned( 8,8)),
			5570 => std_logic_vector(to_unsigned( 30,8)),
			5571 => std_logic_vector(to_unsigned( 76,8)),
			5572 => std_logic_vector(to_unsigned( 81,8)),
			5573 => std_logic_vector(to_unsigned( 30,8)),
			5574 => std_logic_vector(to_unsigned( 134,8)),
			5575 => std_logic_vector(to_unsigned( 43,8)),
			5576 => std_logic_vector(to_unsigned( 58,8)),
			5577 => std_logic_vector(to_unsigned( 12,8)),
			5578 => std_logic_vector(to_unsigned( 242,8)),
			5579 => std_logic_vector(to_unsigned( 120,8)),
			5580 => std_logic_vector(to_unsigned( 79,8)),
			5581 => std_logic_vector(to_unsigned( 103,8)),
			5582 => std_logic_vector(to_unsigned( 140,8)),
			5583 => std_logic_vector(to_unsigned( 143,8)),
			5584 => std_logic_vector(to_unsigned( 219,8)),
			5585 => std_logic_vector(to_unsigned( 125,8)),
			5586 => std_logic_vector(to_unsigned( 190,8)),
			5587 => std_logic_vector(to_unsigned( 203,8)),
			5588 => std_logic_vector(to_unsigned( 79,8)),
			5589 => std_logic_vector(to_unsigned( 236,8)),
			5590 => std_logic_vector(to_unsigned( 237,8)),
			5591 => std_logic_vector(to_unsigned( 107,8)),
			5592 => std_logic_vector(to_unsigned( 98,8)),
			5593 => std_logic_vector(to_unsigned( 63,8)),
			5594 => std_logic_vector(to_unsigned( 238,8)),
			5595 => std_logic_vector(to_unsigned( 244,8)),
			5596 => std_logic_vector(to_unsigned( 64,8)),
			5597 => std_logic_vector(to_unsigned( 119,8)),
			5598 => std_logic_vector(to_unsigned( 81,8)),
			5599 => std_logic_vector(to_unsigned( 103,8)),
			5600 => std_logic_vector(to_unsigned( 215,8)),
			5601 => std_logic_vector(to_unsigned( 194,8)),
			5602 => std_logic_vector(to_unsigned( 223,8)),
			5603 => std_logic_vector(to_unsigned( 12,8)),
			5604 => std_logic_vector(to_unsigned( 212,8)),
			5605 => std_logic_vector(to_unsigned( 223,8)),
			5606 => std_logic_vector(to_unsigned( 244,8)),
			5607 => std_logic_vector(to_unsigned( 229,8)),
			5608 => std_logic_vector(to_unsigned( 31,8)),
			5609 => std_logic_vector(to_unsigned( 80,8)),
			5610 => std_logic_vector(to_unsigned( 151,8)),
			5611 => std_logic_vector(to_unsigned( 120,8)),
			5612 => std_logic_vector(to_unsigned( 56,8)),
			5613 => std_logic_vector(to_unsigned( 241,8)),
			5614 => std_logic_vector(to_unsigned( 156,8)),
			5615 => std_logic_vector(to_unsigned( 196,8)),
			5616 => std_logic_vector(to_unsigned( 225,8)),
			5617 => std_logic_vector(to_unsigned( 199,8)),
			5618 => std_logic_vector(to_unsigned( 166,8)),
			5619 => std_logic_vector(to_unsigned( 220,8)),
			5620 => std_logic_vector(to_unsigned( 154,8)),
			5621 => std_logic_vector(to_unsigned( 99,8)),
			5622 => std_logic_vector(to_unsigned( 73,8)),
			5623 => std_logic_vector(to_unsigned( 212,8)),
			5624 => std_logic_vector(to_unsigned( 109,8)),
			5625 => std_logic_vector(to_unsigned( 106,8)),
			5626 => std_logic_vector(to_unsigned( 194,8)),
			5627 => std_logic_vector(to_unsigned( 16,8)),
			5628 => std_logic_vector(to_unsigned( 43,8)),
			5629 => std_logic_vector(to_unsigned( 55,8)),
			5630 => std_logic_vector(to_unsigned( 176,8)),
			5631 => std_logic_vector(to_unsigned( 22,8)),
			5632 => std_logic_vector(to_unsigned( 61,8)),
			5633 => std_logic_vector(to_unsigned( 99,8)),
			5634 => std_logic_vector(to_unsigned( 27,8)),
			5635 => std_logic_vector(to_unsigned( 162,8)),
			5636 => std_logic_vector(to_unsigned( 205,8)),
			5637 => std_logic_vector(to_unsigned( 158,8)),
			5638 => std_logic_vector(to_unsigned( 217,8)),
			5639 => std_logic_vector(to_unsigned( 63,8)),
			5640 => std_logic_vector(to_unsigned( 156,8)),
			5641 => std_logic_vector(to_unsigned( 16,8)),
			5642 => std_logic_vector(to_unsigned( 135,8)),
			5643 => std_logic_vector(to_unsigned( 83,8)),
			5644 => std_logic_vector(to_unsigned( 149,8)),
			5645 => std_logic_vector(to_unsigned( 196,8)),
			5646 => std_logic_vector(to_unsigned( 171,8)),
			5647 => std_logic_vector(to_unsigned( 175,8)),
			5648 => std_logic_vector(to_unsigned( 190,8)),
			5649 => std_logic_vector(to_unsigned( 29,8)),
			5650 => std_logic_vector(to_unsigned( 54,8)),
			5651 => std_logic_vector(to_unsigned( 86,8)),
			5652 => std_logic_vector(to_unsigned( 230,8)),
			5653 => std_logic_vector(to_unsigned( 132,8)),
			5654 => std_logic_vector(to_unsigned( 39,8)),
			5655 => std_logic_vector(to_unsigned( 109,8)),
			5656 => std_logic_vector(to_unsigned( 194,8)),
			5657 => std_logic_vector(to_unsigned( 72,8)),
			5658 => std_logic_vector(to_unsigned( 206,8)),
			5659 => std_logic_vector(to_unsigned( 157,8)),
			5660 => std_logic_vector(to_unsigned( 80,8)),
			5661 => std_logic_vector(to_unsigned( 144,8)),
			5662 => std_logic_vector(to_unsigned( 125,8)),
			5663 => std_logic_vector(to_unsigned( 114,8)),
			5664 => std_logic_vector(to_unsigned( 5,8)),
			5665 => std_logic_vector(to_unsigned( 230,8)),
			5666 => std_logic_vector(to_unsigned( 61,8)),
			5667 => std_logic_vector(to_unsigned( 246,8)),
			5668 => std_logic_vector(to_unsigned( 72,8)),
			5669 => std_logic_vector(to_unsigned( 13,8)),
			5670 => std_logic_vector(to_unsigned( 87,8)),
			5671 => std_logic_vector(to_unsigned( 58,8)),
			5672 => std_logic_vector(to_unsigned( 65,8)),
			5673 => std_logic_vector(to_unsigned( 152,8)),
			5674 => std_logic_vector(to_unsigned( 247,8)),
			5675 => std_logic_vector(to_unsigned( 183,8)),
			5676 => std_logic_vector(to_unsigned( 105,8)),
			5677 => std_logic_vector(to_unsigned( 104,8)),
			5678 => std_logic_vector(to_unsigned( 96,8)),
			5679 => std_logic_vector(to_unsigned( 197,8)),
			5680 => std_logic_vector(to_unsigned( 35,8)),
			5681 => std_logic_vector(to_unsigned( 20,8)),
			5682 => std_logic_vector(to_unsigned( 192,8)),
			5683 => std_logic_vector(to_unsigned( 173,8)),
			5684 => std_logic_vector(to_unsigned( 250,8)),
			5685 => std_logic_vector(to_unsigned( 253,8)),
			5686 => std_logic_vector(to_unsigned( 60,8)),
			5687 => std_logic_vector(to_unsigned( 227,8)),
			5688 => std_logic_vector(to_unsigned( 74,8)),
			5689 => std_logic_vector(to_unsigned( 172,8)),
			5690 => std_logic_vector(to_unsigned( 139,8)),
			5691 => std_logic_vector(to_unsigned( 190,8)),
			5692 => std_logic_vector(to_unsigned( 50,8)),
			5693 => std_logic_vector(to_unsigned( 60,8)),
			5694 => std_logic_vector(to_unsigned( 12,8)),
			5695 => std_logic_vector(to_unsigned( 253,8)),
			5696 => std_logic_vector(to_unsigned( 122,8)),
			5697 => std_logic_vector(to_unsigned( 121,8)),
			5698 => std_logic_vector(to_unsigned( 228,8)),
			5699 => std_logic_vector(to_unsigned( 133,8)),
			5700 => std_logic_vector(to_unsigned( 141,8)),
			5701 => std_logic_vector(to_unsigned( 89,8)),
			5702 => std_logic_vector(to_unsigned( 43,8)),
			5703 => std_logic_vector(to_unsigned( 189,8)),
			5704 => std_logic_vector(to_unsigned( 236,8)),
			5705 => std_logic_vector(to_unsigned( 125,8)),
			5706 => std_logic_vector(to_unsigned( 57,8)),
			5707 => std_logic_vector(to_unsigned( 8,8)),
			5708 => std_logic_vector(to_unsigned( 247,8)),
			5709 => std_logic_vector(to_unsigned( 24,8)),
			5710 => std_logic_vector(to_unsigned( 124,8)),
			5711 => std_logic_vector(to_unsigned( 214,8)),
			5712 => std_logic_vector(to_unsigned( 130,8)),
			5713 => std_logic_vector(to_unsigned( 177,8)),
			5714 => std_logic_vector(to_unsigned( 202,8)),
			5715 => std_logic_vector(to_unsigned( 66,8)),
			5716 => std_logic_vector(to_unsigned( 68,8)),
			5717 => std_logic_vector(to_unsigned( 153,8)),
			5718 => std_logic_vector(to_unsigned( 252,8)),
			5719 => std_logic_vector(to_unsigned( 13,8)),
			5720 => std_logic_vector(to_unsigned( 25,8)),
			5721 => std_logic_vector(to_unsigned( 94,8)),
			5722 => std_logic_vector(to_unsigned( 125,8)),
			5723 => std_logic_vector(to_unsigned( 202,8)),
			5724 => std_logic_vector(to_unsigned( 88,8)),
			5725 => std_logic_vector(to_unsigned( 149,8)),
			5726 => std_logic_vector(to_unsigned( 103,8)),
			5727 => std_logic_vector(to_unsigned( 138,8)),
			5728 => std_logic_vector(to_unsigned( 64,8)),
			5729 => std_logic_vector(to_unsigned( 67,8)),
			5730 => std_logic_vector(to_unsigned( 214,8)),
			5731 => std_logic_vector(to_unsigned( 235,8)),
			5732 => std_logic_vector(to_unsigned( 189,8)),
			5733 => std_logic_vector(to_unsigned( 52,8)),
			5734 => std_logic_vector(to_unsigned( 70,8)),
			5735 => std_logic_vector(to_unsigned( 191,8)),
			5736 => std_logic_vector(to_unsigned( 104,8)),
			5737 => std_logic_vector(to_unsigned( 202,8)),
			5738 => std_logic_vector(to_unsigned( 205,8)),
			5739 => std_logic_vector(to_unsigned( 54,8)),
			5740 => std_logic_vector(to_unsigned( 180,8)),
			5741 => std_logic_vector(to_unsigned( 168,8)),
			5742 => std_logic_vector(to_unsigned( 192,8)),
			5743 => std_logic_vector(to_unsigned( 89,8)),
			5744 => std_logic_vector(to_unsigned( 58,8)),
			5745 => std_logic_vector(to_unsigned( 10,8)),
			5746 => std_logic_vector(to_unsigned( 217,8)),
			5747 => std_logic_vector(to_unsigned( 32,8)),
			5748 => std_logic_vector(to_unsigned( 147,8)),
			5749 => std_logic_vector(to_unsigned( 26,8)),
			5750 => std_logic_vector(to_unsigned( 124,8)),
			5751 => std_logic_vector(to_unsigned( 134,8)),
			5752 => std_logic_vector(to_unsigned( 224,8)),
			5753 => std_logic_vector(to_unsigned( 76,8)),
			5754 => std_logic_vector(to_unsigned( 161,8)),
			5755 => std_logic_vector(to_unsigned( 122,8)),
			5756 => std_logic_vector(to_unsigned( 202,8)),
			5757 => std_logic_vector(to_unsigned( 56,8)),
			5758 => std_logic_vector(to_unsigned( 25,8)),
			5759 => std_logic_vector(to_unsigned( 77,8)),
			5760 => std_logic_vector(to_unsigned( 118,8)),
			5761 => std_logic_vector(to_unsigned( 156,8)),
			5762 => std_logic_vector(to_unsigned( 107,8)),
			5763 => std_logic_vector(to_unsigned( 30,8)),
			5764 => std_logic_vector(to_unsigned( 195,8)),
			5765 => std_logic_vector(to_unsigned( 116,8)),
			5766 => std_logic_vector(to_unsigned( 188,8)),
			5767 => std_logic_vector(to_unsigned( 219,8)),
			5768 => std_logic_vector(to_unsigned( 248,8)),
			5769 => std_logic_vector(to_unsigned( 109,8)),
			5770 => std_logic_vector(to_unsigned( 219,8)),
			5771 => std_logic_vector(to_unsigned( 127,8)),
			5772 => std_logic_vector(to_unsigned( 105,8)),
			5773 => std_logic_vector(to_unsigned( 215,8)),
			5774 => std_logic_vector(to_unsigned( 69,8)),
			5775 => std_logic_vector(to_unsigned( 124,8)),
			5776 => std_logic_vector(to_unsigned( 123,8)),
			5777 => std_logic_vector(to_unsigned( 133,8)),
			5778 => std_logic_vector(to_unsigned( 125,8)),
			5779 => std_logic_vector(to_unsigned( 156,8)),
			5780 => std_logic_vector(to_unsigned( 62,8)),
			5781 => std_logic_vector(to_unsigned( 145,8)),
			5782 => std_logic_vector(to_unsigned( 53,8)),
			5783 => std_logic_vector(to_unsigned( 11,8)),
			5784 => std_logic_vector(to_unsigned( 31,8)),
			5785 => std_logic_vector(to_unsigned( 86,8)),
			5786 => std_logic_vector(to_unsigned( 137,8)),
			5787 => std_logic_vector(to_unsigned( 39,8)),
			5788 => std_logic_vector(to_unsigned( 176,8)),
			5789 => std_logic_vector(to_unsigned( 167,8)),
			5790 => std_logic_vector(to_unsigned( 92,8)),
			5791 => std_logic_vector(to_unsigned( 120,8)),
			5792 => std_logic_vector(to_unsigned( 49,8)),
			5793 => std_logic_vector(to_unsigned( 243,8)),
			5794 => std_logic_vector(to_unsigned( 255,8)),
			5795 => std_logic_vector(to_unsigned( 25,8)),
			5796 => std_logic_vector(to_unsigned( 231,8)),
			5797 => std_logic_vector(to_unsigned( 240,8)),
			5798 => std_logic_vector(to_unsigned( 254,8)),
			5799 => std_logic_vector(to_unsigned( 243,8)),
			5800 => std_logic_vector(to_unsigned( 134,8)),
			5801 => std_logic_vector(to_unsigned( 135,8)),
			5802 => std_logic_vector(to_unsigned( 96,8)),
			5803 => std_logic_vector(to_unsigned( 22,8)),
			5804 => std_logic_vector(to_unsigned( 8,8)),
			5805 => std_logic_vector(to_unsigned( 216,8)),
			5806 => std_logic_vector(to_unsigned( 87,8)),
			5807 => std_logic_vector(to_unsigned( 57,8)),
			5808 => std_logic_vector(to_unsigned( 137,8)),
			5809 => std_logic_vector(to_unsigned( 150,8)),
			5810 => std_logic_vector(to_unsigned( 68,8)),
			5811 => std_logic_vector(to_unsigned( 74,8)),
			5812 => std_logic_vector(to_unsigned( 141,8)),
			5813 => std_logic_vector(to_unsigned( 233,8)),
			5814 => std_logic_vector(to_unsigned( 4,8)),
			5815 => std_logic_vector(to_unsigned( 42,8)),
			5816 => std_logic_vector(to_unsigned( 83,8)),
			5817 => std_logic_vector(to_unsigned( 220,8)),
			5818 => std_logic_vector(to_unsigned( 201,8)),
			5819 => std_logic_vector(to_unsigned( 56,8)),
			5820 => std_logic_vector(to_unsigned( 219,8)),
			5821 => std_logic_vector(to_unsigned( 78,8)),
			5822 => std_logic_vector(to_unsigned( 239,8)),
			5823 => std_logic_vector(to_unsigned( 148,8)),
			5824 => std_logic_vector(to_unsigned( 136,8)),
			5825 => std_logic_vector(to_unsigned( 186,8)),
			5826 => std_logic_vector(to_unsigned( 52,8)),
			5827 => std_logic_vector(to_unsigned( 40,8)),
			5828 => std_logic_vector(to_unsigned( 29,8)),
			5829 => std_logic_vector(to_unsigned( 173,8)),
			5830 => std_logic_vector(to_unsigned( 119,8)),
			5831 => std_logic_vector(to_unsigned( 11,8)),
			5832 => std_logic_vector(to_unsigned( 231,8)),
			5833 => std_logic_vector(to_unsigned( 26,8)),
			5834 => std_logic_vector(to_unsigned( 23,8)),
			5835 => std_logic_vector(to_unsigned( 55,8)),
			5836 => std_logic_vector(to_unsigned( 121,8)),
			5837 => std_logic_vector(to_unsigned( 141,8)),
			5838 => std_logic_vector(to_unsigned( 34,8)),
			5839 => std_logic_vector(to_unsigned( 42,8)),
			5840 => std_logic_vector(to_unsigned( 141,8)),
			5841 => std_logic_vector(to_unsigned( 113,8)),
			5842 => std_logic_vector(to_unsigned( 198,8)),
			5843 => std_logic_vector(to_unsigned( 51,8)),
			5844 => std_logic_vector(to_unsigned( 209,8)),
			5845 => std_logic_vector(to_unsigned( 181,8)),
			5846 => std_logic_vector(to_unsigned( 91,8)),
			5847 => std_logic_vector(to_unsigned( 224,8)),
			5848 => std_logic_vector(to_unsigned( 34,8)),
			5849 => std_logic_vector(to_unsigned( 183,8)),
			5850 => std_logic_vector(to_unsigned( 63,8)),
			5851 => std_logic_vector(to_unsigned( 47,8)),
			5852 => std_logic_vector(to_unsigned( 70,8)),
			5853 => std_logic_vector(to_unsigned( 119,8)),
			5854 => std_logic_vector(to_unsigned( 17,8)),
			5855 => std_logic_vector(to_unsigned( 243,8)),
			5856 => std_logic_vector(to_unsigned( 210,8)),
			5857 => std_logic_vector(to_unsigned( 163,8)),
			5858 => std_logic_vector(to_unsigned( 179,8)),
			5859 => std_logic_vector(to_unsigned( 168,8)),
			5860 => std_logic_vector(to_unsigned( 208,8)),
			5861 => std_logic_vector(to_unsigned( 192,8)),
			5862 => std_logic_vector(to_unsigned( 222,8)),
			5863 => std_logic_vector(to_unsigned( 87,8)),
			5864 => std_logic_vector(to_unsigned( 113,8)),
			5865 => std_logic_vector(to_unsigned( 132,8)),
			5866 => std_logic_vector(to_unsigned( 17,8)),
			5867 => std_logic_vector(to_unsigned( 62,8)),
			5868 => std_logic_vector(to_unsigned( 23,8)),
			5869 => std_logic_vector(to_unsigned( 198,8)),
			5870 => std_logic_vector(to_unsigned( 19,8)),
			5871 => std_logic_vector(to_unsigned( 152,8)),
			5872 => std_logic_vector(to_unsigned( 14,8)),
			5873 => std_logic_vector(to_unsigned( 170,8)),
			5874 => std_logic_vector(to_unsigned( 124,8)),
			5875 => std_logic_vector(to_unsigned( 24,8)),
			5876 => std_logic_vector(to_unsigned( 169,8)),
			5877 => std_logic_vector(to_unsigned( 38,8)),
			5878 => std_logic_vector(to_unsigned( 168,8)),
			5879 => std_logic_vector(to_unsigned( 134,8)),
			5880 => std_logic_vector(to_unsigned( 116,8)),
			5881 => std_logic_vector(to_unsigned( 89,8)),
			5882 => std_logic_vector(to_unsigned( 33,8)),
			5883 => std_logic_vector(to_unsigned( 208,8)),
			5884 => std_logic_vector(to_unsigned( 188,8)),
			5885 => std_logic_vector(to_unsigned( 130,8)),
			5886 => std_logic_vector(to_unsigned( 127,8)),
			5887 => std_logic_vector(to_unsigned( 173,8)),
			5888 => std_logic_vector(to_unsigned( 142,8)),
			5889 => std_logic_vector(to_unsigned( 205,8)),
			5890 => std_logic_vector(to_unsigned( 3,8)),
			5891 => std_logic_vector(to_unsigned( 208,8)),
			5892 => std_logic_vector(to_unsigned( 126,8)),
			5893 => std_logic_vector(to_unsigned( 72,8)),
			5894 => std_logic_vector(to_unsigned( 191,8)),
			5895 => std_logic_vector(to_unsigned( 139,8)),
			5896 => std_logic_vector(to_unsigned( 209,8)),
			5897 => std_logic_vector(to_unsigned( 175,8)),
			5898 => std_logic_vector(to_unsigned( 89,8)),
			5899 => std_logic_vector(to_unsigned( 182,8)),
			5900 => std_logic_vector(to_unsigned( 123,8)),
			5901 => std_logic_vector(to_unsigned( 113,8)),
			5902 => std_logic_vector(to_unsigned( 239,8)),
			5903 => std_logic_vector(to_unsigned( 156,8)),
			5904 => std_logic_vector(to_unsigned( 252,8)),
			5905 => std_logic_vector(to_unsigned( 228,8)),
			5906 => std_logic_vector(to_unsigned( 252,8)),
			5907 => std_logic_vector(to_unsigned( 191,8)),
			5908 => std_logic_vector(to_unsigned( 4,8)),
			5909 => std_logic_vector(to_unsigned( 69,8)),
			5910 => std_logic_vector(to_unsigned( 28,8)),
			5911 => std_logic_vector(to_unsigned( 39,8)),
			5912 => std_logic_vector(to_unsigned( 162,8)),
			5913 => std_logic_vector(to_unsigned( 110,8)),
			5914 => std_logic_vector(to_unsigned( 152,8)),
			5915 => std_logic_vector(to_unsigned( 178,8)),
			5916 => std_logic_vector(to_unsigned( 122,8)),
			5917 => std_logic_vector(to_unsigned( 99,8)),
			5918 => std_logic_vector(to_unsigned( 140,8)),
			5919 => std_logic_vector(to_unsigned( 33,8)),
			5920 => std_logic_vector(to_unsigned( 214,8)),
			5921 => std_logic_vector(to_unsigned( 116,8)),
			5922 => std_logic_vector(to_unsigned( 73,8)),
			5923 => std_logic_vector(to_unsigned( 133,8)),
			5924 => std_logic_vector(to_unsigned( 133,8)),
			5925 => std_logic_vector(to_unsigned( 56,8)),
			5926 => std_logic_vector(to_unsigned( 30,8)),
			5927 => std_logic_vector(to_unsigned( 140,8)),
			5928 => std_logic_vector(to_unsigned( 245,8)),
			5929 => std_logic_vector(to_unsigned( 195,8)),
			5930 => std_logic_vector(to_unsigned( 116,8)),
			5931 => std_logic_vector(to_unsigned( 11,8)),
			5932 => std_logic_vector(to_unsigned( 130,8)),
			5933 => std_logic_vector(to_unsigned( 179,8)),
			5934 => std_logic_vector(to_unsigned( 109,8)),
			5935 => std_logic_vector(to_unsigned( 51,8)),
			5936 => std_logic_vector(to_unsigned( 251,8)),
			5937 => std_logic_vector(to_unsigned( 21,8)),
			5938 => std_logic_vector(to_unsigned( 41,8)),
			5939 => std_logic_vector(to_unsigned( 89,8)),
			5940 => std_logic_vector(to_unsigned( 34,8)),
			5941 => std_logic_vector(to_unsigned( 243,8)),
			5942 => std_logic_vector(to_unsigned( 44,8)),
			5943 => std_logic_vector(to_unsigned( 136,8)),
			5944 => std_logic_vector(to_unsigned( 130,8)),
			5945 => std_logic_vector(to_unsigned( 110,8)),
			5946 => std_logic_vector(to_unsigned( 247,8)),
			5947 => std_logic_vector(to_unsigned( 14,8)),
			5948 => std_logic_vector(to_unsigned( 203,8)),
			5949 => std_logic_vector(to_unsigned( 61,8)),
			5950 => std_logic_vector(to_unsigned( 93,8)),
			5951 => std_logic_vector(to_unsigned( 184,8)),
			5952 => std_logic_vector(to_unsigned( 53,8)),
			5953 => std_logic_vector(to_unsigned( 127,8)),
			5954 => std_logic_vector(to_unsigned( 192,8)),
			5955 => std_logic_vector(to_unsigned( 164,8)),
			5956 => std_logic_vector(to_unsigned( 60,8)),
			5957 => std_logic_vector(to_unsigned( 142,8)),
			5958 => std_logic_vector(to_unsigned( 122,8)),
			5959 => std_logic_vector(to_unsigned( 108,8)),
			5960 => std_logic_vector(to_unsigned( 245,8)),
			5961 => std_logic_vector(to_unsigned( 83,8)),
			5962 => std_logic_vector(to_unsigned( 128,8)),
			5963 => std_logic_vector(to_unsigned( 45,8)),
			5964 => std_logic_vector(to_unsigned( 31,8)),
			5965 => std_logic_vector(to_unsigned( 194,8)),
			5966 => std_logic_vector(to_unsigned( 106,8)),
			5967 => std_logic_vector(to_unsigned( 112,8)),
			5968 => std_logic_vector(to_unsigned( 172,8)),
			5969 => std_logic_vector(to_unsigned( 130,8)),
			5970 => std_logic_vector(to_unsigned( 68,8)),
			5971 => std_logic_vector(to_unsigned( 208,8)),
			5972 => std_logic_vector(to_unsigned( 47,8)),
			5973 => std_logic_vector(to_unsigned( 153,8)),
			5974 => std_logic_vector(to_unsigned( 53,8)),
			5975 => std_logic_vector(to_unsigned( 68,8)),
			5976 => std_logic_vector(to_unsigned( 246,8)),
			5977 => std_logic_vector(to_unsigned( 119,8)),
			5978 => std_logic_vector(to_unsigned( 63,8)),
			5979 => std_logic_vector(to_unsigned( 168,8)),
			5980 => std_logic_vector(to_unsigned( 242,8)),
			5981 => std_logic_vector(to_unsigned( 161,8)),
			5982 => std_logic_vector(to_unsigned( 118,8)),
			5983 => std_logic_vector(to_unsigned( 40,8)),
			5984 => std_logic_vector(to_unsigned( 96,8)),
			5985 => std_logic_vector(to_unsigned( 210,8)),
			5986 => std_logic_vector(to_unsigned( 92,8)),
			5987 => std_logic_vector(to_unsigned( 17,8)),
			5988 => std_logic_vector(to_unsigned( 234,8)),
			5989 => std_logic_vector(to_unsigned( 17,8)),
			5990 => std_logic_vector(to_unsigned( 230,8)),
			5991 => std_logic_vector(to_unsigned( 8,8)),
			5992 => std_logic_vector(to_unsigned( 236,8)),
			5993 => std_logic_vector(to_unsigned( 114,8)),
			5994 => std_logic_vector(to_unsigned( 17,8)),
			5995 => std_logic_vector(to_unsigned( 168,8)),
			5996 => std_logic_vector(to_unsigned( 149,8)),
			5997 => std_logic_vector(to_unsigned( 75,8)),
			5998 => std_logic_vector(to_unsigned( 86,8)),
			5999 => std_logic_vector(to_unsigned( 234,8)),
			6000 => std_logic_vector(to_unsigned( 9,8)),
			6001 => std_logic_vector(to_unsigned( 228,8)),
			6002 => std_logic_vector(to_unsigned( 25,8)),
			6003 => std_logic_vector(to_unsigned( 2,8)),
			6004 => std_logic_vector(to_unsigned( 61,8)),
			6005 => std_logic_vector(to_unsigned( 54,8)),
			6006 => std_logic_vector(to_unsigned( 121,8)),
			6007 => std_logic_vector(to_unsigned( 27,8)),
			6008 => std_logic_vector(to_unsigned( 142,8)),
			6009 => std_logic_vector(to_unsigned( 87,8)),
			6010 => std_logic_vector(to_unsigned( 117,8)),
			6011 => std_logic_vector(to_unsigned( 56,8)),
			6012 => std_logic_vector(to_unsigned( 249,8)),
			6013 => std_logic_vector(to_unsigned( 241,8)),
			6014 => std_logic_vector(to_unsigned( 107,8)),
			6015 => std_logic_vector(to_unsigned( 143,8)),
			6016 => std_logic_vector(to_unsigned( 184,8)),
			6017 => std_logic_vector(to_unsigned( 1,8)),
			6018 => std_logic_vector(to_unsigned( 106,8)),
			6019 => std_logic_vector(to_unsigned( 185,8)),
			6020 => std_logic_vector(to_unsigned( 78,8)),
			6021 => std_logic_vector(to_unsigned( 86,8)),
			6022 => std_logic_vector(to_unsigned( 145,8)),
			6023 => std_logic_vector(to_unsigned( 212,8)),
			6024 => std_logic_vector(to_unsigned( 59,8)),
			6025 => std_logic_vector(to_unsigned( 74,8)),
			6026 => std_logic_vector(to_unsigned( 235,8)),
			6027 => std_logic_vector(to_unsigned( 208,8)),
			6028 => std_logic_vector(to_unsigned( 98,8)),
			6029 => std_logic_vector(to_unsigned( 235,8)),
			6030 => std_logic_vector(to_unsigned( 52,8)),
			6031 => std_logic_vector(to_unsigned( 221,8)),
			6032 => std_logic_vector(to_unsigned( 196,8)),
			6033 => std_logic_vector(to_unsigned( 200,8)),
			6034 => std_logic_vector(to_unsigned( 171,8)),
			6035 => std_logic_vector(to_unsigned( 96,8)),
			6036 => std_logic_vector(to_unsigned( 252,8)),
			6037 => std_logic_vector(to_unsigned( 50,8)),
			6038 => std_logic_vector(to_unsigned( 159,8)),
			6039 => std_logic_vector(to_unsigned( 197,8)),
			6040 => std_logic_vector(to_unsigned( 71,8)),
			6041 => std_logic_vector(to_unsigned( 108,8)),
			6042 => std_logic_vector(to_unsigned( 215,8)),
			6043 => std_logic_vector(to_unsigned( 51,8)),
			6044 => std_logic_vector(to_unsigned( 143,8)),
			6045 => std_logic_vector(to_unsigned( 250,8)),
			6046 => std_logic_vector(to_unsigned( 32,8)),
			6047 => std_logic_vector(to_unsigned( 22,8)),
			6048 => std_logic_vector(to_unsigned( 177,8)),
			6049 => std_logic_vector(to_unsigned( 130,8)),
			6050 => std_logic_vector(to_unsigned( 113,8)),
			6051 => std_logic_vector(to_unsigned( 70,8)),
			6052 => std_logic_vector(to_unsigned( 255,8)),
			6053 => std_logic_vector(to_unsigned( 23,8)),
			6054 => std_logic_vector(to_unsigned( 190,8)),
			6055 => std_logic_vector(to_unsigned( 210,8)),
			6056 => std_logic_vector(to_unsigned( 101,8)),
			6057 => std_logic_vector(to_unsigned( 72,8)),
			6058 => std_logic_vector(to_unsigned( 68,8)),
			6059 => std_logic_vector(to_unsigned( 189,8)),
			6060 => std_logic_vector(to_unsigned( 27,8)),
			6061 => std_logic_vector(to_unsigned( 239,8)),
			6062 => std_logic_vector(to_unsigned( 91,8)),
			6063 => std_logic_vector(to_unsigned( 157,8)),
			6064 => std_logic_vector(to_unsigned( 29,8)),
			6065 => std_logic_vector(to_unsigned( 206,8)),
			6066 => std_logic_vector(to_unsigned( 51,8)),
			6067 => std_logic_vector(to_unsigned( 47,8)),
			6068 => std_logic_vector(to_unsigned( 186,8)),
			6069 => std_logic_vector(to_unsigned( 167,8)),
			6070 => std_logic_vector(to_unsigned( 197,8)),
			6071 => std_logic_vector(to_unsigned( 206,8)),
			6072 => std_logic_vector(to_unsigned( 161,8)),
			6073 => std_logic_vector(to_unsigned( 197,8)),
			6074 => std_logic_vector(to_unsigned( 19,8)),
			6075 => std_logic_vector(to_unsigned( 217,8)),
			6076 => std_logic_vector(to_unsigned( 113,8)),
			6077 => std_logic_vector(to_unsigned( 240,8)),
			6078 => std_logic_vector(to_unsigned( 208,8)),
			6079 => std_logic_vector(to_unsigned( 158,8)),
			6080 => std_logic_vector(to_unsigned( 95,8)),
			6081 => std_logic_vector(to_unsigned( 74,8)),
			6082 => std_logic_vector(to_unsigned( 223,8)),
			6083 => std_logic_vector(to_unsigned( 10,8)),
			6084 => std_logic_vector(to_unsigned( 116,8)),
			6085 => std_logic_vector(to_unsigned( 181,8)),
			6086 => std_logic_vector(to_unsigned( 167,8)),
			6087 => std_logic_vector(to_unsigned( 71,8)),
			6088 => std_logic_vector(to_unsigned( 175,8)),
			6089 => std_logic_vector(to_unsigned( 45,8)),
			6090 => std_logic_vector(to_unsigned( 215,8)),
			6091 => std_logic_vector(to_unsigned( 186,8)),
			6092 => std_logic_vector(to_unsigned( 107,8)),
			6093 => std_logic_vector(to_unsigned( 161,8)),
			6094 => std_logic_vector(to_unsigned( 225,8)),
			6095 => std_logic_vector(to_unsigned( 72,8)),
			6096 => std_logic_vector(to_unsigned( 23,8)),
			6097 => std_logic_vector(to_unsigned( 91,8)),
			6098 => std_logic_vector(to_unsigned( 152,8)),
			6099 => std_logic_vector(to_unsigned( 195,8)),
			6100 => std_logic_vector(to_unsigned( 105,8)),
			6101 => std_logic_vector(to_unsigned( 196,8)),
			6102 => std_logic_vector(to_unsigned( 204,8)),
			6103 => std_logic_vector(to_unsigned( 11,8)),
			6104 => std_logic_vector(to_unsigned( 224,8)),
			6105 => std_logic_vector(to_unsigned( 152,8)),
			6106 => std_logic_vector(to_unsigned( 25,8)),
			6107 => std_logic_vector(to_unsigned( 71,8)),
			6108 => std_logic_vector(to_unsigned( 254,8)),
			6109 => std_logic_vector(to_unsigned( 31,8)),
			6110 => std_logic_vector(to_unsigned( 207,8)),
			6111 => std_logic_vector(to_unsigned( 190,8)),
			6112 => std_logic_vector(to_unsigned( 105,8)),
			6113 => std_logic_vector(to_unsigned( 79,8)),
			6114 => std_logic_vector(to_unsigned( 180,8)),
			6115 => std_logic_vector(to_unsigned( 157,8)),
			6116 => std_logic_vector(to_unsigned( 168,8)),
			6117 => std_logic_vector(to_unsigned( 156,8)),
			6118 => std_logic_vector(to_unsigned( 48,8)),
			6119 => std_logic_vector(to_unsigned( 3,8)),
			6120 => std_logic_vector(to_unsigned( 58,8)),
			6121 => std_logic_vector(to_unsigned( 114,8)),
			6122 => std_logic_vector(to_unsigned( 48,8)),
			6123 => std_logic_vector(to_unsigned( 212,8)),
			6124 => std_logic_vector(to_unsigned( 0,8)),
			6125 => std_logic_vector(to_unsigned( 189,8)),
			6126 => std_logic_vector(to_unsigned( 93,8)),
			6127 => std_logic_vector(to_unsigned( 53,8)),
			6128 => std_logic_vector(to_unsigned( 219,8)),
			6129 => std_logic_vector(to_unsigned( 224,8)),
			6130 => std_logic_vector(to_unsigned( 247,8)),
			6131 => std_logic_vector(to_unsigned( 105,8)),
			6132 => std_logic_vector(to_unsigned( 240,8)),
			6133 => std_logic_vector(to_unsigned( 208,8)),
			6134 => std_logic_vector(to_unsigned( 15,8)),
			6135 => std_logic_vector(to_unsigned( 254,8)),
			6136 => std_logic_vector(to_unsigned( 211,8)),
			6137 => std_logic_vector(to_unsigned( 200,8)),
			6138 => std_logic_vector(to_unsigned( 244,8)),
			6139 => std_logic_vector(to_unsigned( 5,8)),
			6140 => std_logic_vector(to_unsigned( 63,8)),
			6141 => std_logic_vector(to_unsigned( 27,8)),
			6142 => std_logic_vector(to_unsigned( 149,8)),
			6143 => std_logic_vector(to_unsigned( 173,8)),
			6144 => std_logic_vector(to_unsigned( 45,8)),
			6145 => std_logic_vector(to_unsigned( 223,8)),
			6146 => std_logic_vector(to_unsigned( 136,8)),
			6147 => std_logic_vector(to_unsigned( 67,8)),
			6148 => std_logic_vector(to_unsigned( 225,8)),
			6149 => std_logic_vector(to_unsigned( 213,8)),
			6150 => std_logic_vector(to_unsigned( 40,8)),
			6151 => std_logic_vector(to_unsigned( 65,8)),
			6152 => std_logic_vector(to_unsigned( 248,8)),
			6153 => std_logic_vector(to_unsigned( 91,8)),
			6154 => std_logic_vector(to_unsigned( 178,8)),
			6155 => std_logic_vector(to_unsigned( 15,8)),
			6156 => std_logic_vector(to_unsigned( 193,8)),
			6157 => std_logic_vector(to_unsigned( 105,8)),
			6158 => std_logic_vector(to_unsigned( 248,8)),
			6159 => std_logic_vector(to_unsigned( 129,8)),
			6160 => std_logic_vector(to_unsigned( 142,8)),
			6161 => std_logic_vector(to_unsigned( 50,8)),
			6162 => std_logic_vector(to_unsigned( 111,8)),
			6163 => std_logic_vector(to_unsigned( 173,8)),
			6164 => std_logic_vector(to_unsigned( 158,8)),
			6165 => std_logic_vector(to_unsigned( 87,8)),
			6166 => std_logic_vector(to_unsigned( 226,8)),
			6167 => std_logic_vector(to_unsigned( 204,8)),
			6168 => std_logic_vector(to_unsigned( 47,8)),
			6169 => std_logic_vector(to_unsigned( 104,8)),
			6170 => std_logic_vector(to_unsigned( 18,8)),
			6171 => std_logic_vector(to_unsigned( 50,8)),
			6172 => std_logic_vector(to_unsigned( 161,8)),
			6173 => std_logic_vector(to_unsigned( 82,8)),
			6174 => std_logic_vector(to_unsigned( 249,8)),
			6175 => std_logic_vector(to_unsigned( 138,8)),
			6176 => std_logic_vector(to_unsigned( 167,8)),
			6177 => std_logic_vector(to_unsigned( 73,8)),
			6178 => std_logic_vector(to_unsigned( 116,8)),
			6179 => std_logic_vector(to_unsigned( 8,8)),
			6180 => std_logic_vector(to_unsigned( 38,8)),
			6181 => std_logic_vector(to_unsigned( 47,8)),
			6182 => std_logic_vector(to_unsigned( 242,8)),
			6183 => std_logic_vector(to_unsigned( 224,8)),
			6184 => std_logic_vector(to_unsigned( 90,8)),
			6185 => std_logic_vector(to_unsigned( 41,8)),
			6186 => std_logic_vector(to_unsigned( 4,8)),
			6187 => std_logic_vector(to_unsigned( 154,8)),
			6188 => std_logic_vector(to_unsigned( 178,8)),
			6189 => std_logic_vector(to_unsigned( 86,8)),
			6190 => std_logic_vector(to_unsigned( 30,8)),
			6191 => std_logic_vector(to_unsigned( 60,8)),
			6192 => std_logic_vector(to_unsigned( 198,8)),
			6193 => std_logic_vector(to_unsigned( 181,8)),
			6194 => std_logic_vector(to_unsigned( 63,8)),
			6195 => std_logic_vector(to_unsigned( 127,8)),
			6196 => std_logic_vector(to_unsigned( 195,8)),
			6197 => std_logic_vector(to_unsigned( 179,8)),
			6198 => std_logic_vector(to_unsigned( 164,8)),
			6199 => std_logic_vector(to_unsigned( 176,8)),
			6200 => std_logic_vector(to_unsigned( 192,8)),
			6201 => std_logic_vector(to_unsigned( 24,8)),
			6202 => std_logic_vector(to_unsigned( 230,8)),
			6203 => std_logic_vector(to_unsigned( 100,8)),
			6204 => std_logic_vector(to_unsigned( 68,8)),
			6205 => std_logic_vector(to_unsigned( 187,8)),
			6206 => std_logic_vector(to_unsigned( 205,8)),
			6207 => std_logic_vector(to_unsigned( 216,8)),
			6208 => std_logic_vector(to_unsigned( 173,8)),
			6209 => std_logic_vector(to_unsigned( 106,8)),
			6210 => std_logic_vector(to_unsigned( 122,8)),
			6211 => std_logic_vector(to_unsigned( 17,8)),
			6212 => std_logic_vector(to_unsigned( 50,8)),
			6213 => std_logic_vector(to_unsigned( 223,8)),
			6214 => std_logic_vector(to_unsigned( 149,8)),
			6215 => std_logic_vector(to_unsigned( 254,8)),
			6216 => std_logic_vector(to_unsigned( 63,8)),
			6217 => std_logic_vector(to_unsigned( 225,8)),
			6218 => std_logic_vector(to_unsigned( 240,8)),
			6219 => std_logic_vector(to_unsigned( 81,8)),
			6220 => std_logic_vector(to_unsigned( 157,8)),
			6221 => std_logic_vector(to_unsigned( 71,8)),
			6222 => std_logic_vector(to_unsigned( 73,8)),
			6223 => std_logic_vector(to_unsigned( 94,8)),
			6224 => std_logic_vector(to_unsigned( 252,8)),
			6225 => std_logic_vector(to_unsigned( 39,8)),
			6226 => std_logic_vector(to_unsigned( 86,8)),
			6227 => std_logic_vector(to_unsigned( 106,8)),
			6228 => std_logic_vector(to_unsigned( 81,8)),
			6229 => std_logic_vector(to_unsigned( 1,8)),
			6230 => std_logic_vector(to_unsigned( 144,8)),
			6231 => std_logic_vector(to_unsigned( 217,8)),
			6232 => std_logic_vector(to_unsigned( 45,8)),
			6233 => std_logic_vector(to_unsigned( 92,8)),
			6234 => std_logic_vector(to_unsigned( 222,8)),
			6235 => std_logic_vector(to_unsigned( 87,8)),
			6236 => std_logic_vector(to_unsigned( 50,8)),
			6237 => std_logic_vector(to_unsigned( 72,8)),
			6238 => std_logic_vector(to_unsigned( 19,8)),
			6239 => std_logic_vector(to_unsigned( 190,8)),
			6240 => std_logic_vector(to_unsigned( 242,8)),
			6241 => std_logic_vector(to_unsigned( 191,8)),
			6242 => std_logic_vector(to_unsigned( 75,8)),
			6243 => std_logic_vector(to_unsigned( 118,8)),
			6244 => std_logic_vector(to_unsigned( 126,8)),
			6245 => std_logic_vector(to_unsigned( 145,8)),
			6246 => std_logic_vector(to_unsigned( 89,8)),
			6247 => std_logic_vector(to_unsigned( 7,8)),
			6248 => std_logic_vector(to_unsigned( 164,8)),
			6249 => std_logic_vector(to_unsigned( 228,8)),
			6250 => std_logic_vector(to_unsigned( 219,8)),
			6251 => std_logic_vector(to_unsigned( 31,8)),
			6252 => std_logic_vector(to_unsigned( 5,8)),
			6253 => std_logic_vector(to_unsigned( 22,8)),
			6254 => std_logic_vector(to_unsigned( 199,8)),
			6255 => std_logic_vector(to_unsigned( 159,8)),
			6256 => std_logic_vector(to_unsigned( 174,8)),
			6257 => std_logic_vector(to_unsigned( 156,8)),
			6258 => std_logic_vector(to_unsigned( 6,8)),
			6259 => std_logic_vector(to_unsigned( 193,8)),
			6260 => std_logic_vector(to_unsigned( 25,8)),
			6261 => std_logic_vector(to_unsigned( 50,8)),
			6262 => std_logic_vector(to_unsigned( 13,8)),
			6263 => std_logic_vector(to_unsigned( 99,8)),
			6264 => std_logic_vector(to_unsigned( 252,8)),
			6265 => std_logic_vector(to_unsigned( 46,8)),
			6266 => std_logic_vector(to_unsigned( 213,8)),
			6267 => std_logic_vector(to_unsigned( 91,8)),
			6268 => std_logic_vector(to_unsigned( 229,8)),
			6269 => std_logic_vector(to_unsigned( 46,8)),
			6270 => std_logic_vector(to_unsigned( 188,8)),
			6271 => std_logic_vector(to_unsigned( 18,8)),
			6272 => std_logic_vector(to_unsigned( 231,8)),
			6273 => std_logic_vector(to_unsigned( 173,8)),
			6274 => std_logic_vector(to_unsigned( 106,8)),
			6275 => std_logic_vector(to_unsigned( 125,8)),
			6276 => std_logic_vector(to_unsigned( 132,8)),
			6277 => std_logic_vector(to_unsigned( 90,8)),
			6278 => std_logic_vector(to_unsigned( 217,8)),
			6279 => std_logic_vector(to_unsigned( 186,8)),
			6280 => std_logic_vector(to_unsigned( 83,8)),
			6281 => std_logic_vector(to_unsigned( 30,8)),
			6282 => std_logic_vector(to_unsigned( 154,8)),
			6283 => std_logic_vector(to_unsigned( 125,8)),
			6284 => std_logic_vector(to_unsigned( 222,8)),
			6285 => std_logic_vector(to_unsigned( 99,8)),
			6286 => std_logic_vector(to_unsigned( 60,8)),
			6287 => std_logic_vector(to_unsigned( 2,8)),
			6288 => std_logic_vector(to_unsigned( 39,8)),
			6289 => std_logic_vector(to_unsigned( 233,8)),
			6290 => std_logic_vector(to_unsigned( 44,8)),
			6291 => std_logic_vector(to_unsigned( 211,8)),
			6292 => std_logic_vector(to_unsigned( 209,8)),
			6293 => std_logic_vector(to_unsigned( 51,8)),
			6294 => std_logic_vector(to_unsigned( 163,8)),
			6295 => std_logic_vector(to_unsigned( 244,8)),
			6296 => std_logic_vector(to_unsigned( 116,8)),
			6297 => std_logic_vector(to_unsigned( 93,8)),
			6298 => std_logic_vector(to_unsigned( 179,8)),
			6299 => std_logic_vector(to_unsigned( 106,8)),
			6300 => std_logic_vector(to_unsigned( 46,8)),
			6301 => std_logic_vector(to_unsigned( 27,8)),
			6302 => std_logic_vector(to_unsigned( 2,8)),
			6303 => std_logic_vector(to_unsigned( 106,8)),
			6304 => std_logic_vector(to_unsigned( 102,8)),
			6305 => std_logic_vector(to_unsigned( 202,8)),
			6306 => std_logic_vector(to_unsigned( 129,8)),
			6307 => std_logic_vector(to_unsigned( 77,8)),
			6308 => std_logic_vector(to_unsigned( 51,8)),
			6309 => std_logic_vector(to_unsigned( 194,8)),
			6310 => std_logic_vector(to_unsigned( 135,8)),
			6311 => std_logic_vector(to_unsigned( 126,8)),
			6312 => std_logic_vector(to_unsigned( 102,8)),
			6313 => std_logic_vector(to_unsigned( 208,8)),
			6314 => std_logic_vector(to_unsigned( 188,8)),
			6315 => std_logic_vector(to_unsigned( 244,8)),
			6316 => std_logic_vector(to_unsigned( 60,8)),
			6317 => std_logic_vector(to_unsigned( 32,8)),
			6318 => std_logic_vector(to_unsigned( 155,8)),
			6319 => std_logic_vector(to_unsigned( 162,8)),
			6320 => std_logic_vector(to_unsigned( 151,8)),
			6321 => std_logic_vector(to_unsigned( 22,8)),
			6322 => std_logic_vector(to_unsigned( 134,8)),
			6323 => std_logic_vector(to_unsigned( 68,8)),
			6324 => std_logic_vector(to_unsigned( 170,8)),
			6325 => std_logic_vector(to_unsigned( 35,8)),
			6326 => std_logic_vector(to_unsigned( 103,8)),
			6327 => std_logic_vector(to_unsigned( 108,8)),
			6328 => std_logic_vector(to_unsigned( 4,8)),
			6329 => std_logic_vector(to_unsigned( 100,8)),
			6330 => std_logic_vector(to_unsigned( 93,8)),
			6331 => std_logic_vector(to_unsigned( 188,8)),
			6332 => std_logic_vector(to_unsigned( 82,8)),
			6333 => std_logic_vector(to_unsigned( 197,8)),
			6334 => std_logic_vector(to_unsigned( 190,8)),
			6335 => std_logic_vector(to_unsigned( 87,8)),
			6336 => std_logic_vector(to_unsigned( 36,8)),
			6337 => std_logic_vector(to_unsigned( 197,8)),
			6338 => std_logic_vector(to_unsigned( 79,8)),
			6339 => std_logic_vector(to_unsigned( 121,8)),
			6340 => std_logic_vector(to_unsigned( 84,8)),
			6341 => std_logic_vector(to_unsigned( 147,8)),
			6342 => std_logic_vector(to_unsigned( 169,8)),
			6343 => std_logic_vector(to_unsigned( 78,8)),
			6344 => std_logic_vector(to_unsigned( 248,8)),
			6345 => std_logic_vector(to_unsigned( 221,8)),
			6346 => std_logic_vector(to_unsigned( 245,8)),
			6347 => std_logic_vector(to_unsigned( 97,8)),
			6348 => std_logic_vector(to_unsigned( 44,8)),
			6349 => std_logic_vector(to_unsigned( 16,8)),
			6350 => std_logic_vector(to_unsigned( 25,8)),
			6351 => std_logic_vector(to_unsigned( 135,8)),
			6352 => std_logic_vector(to_unsigned( 86,8)),
			6353 => std_logic_vector(to_unsigned( 16,8)),
			6354 => std_logic_vector(to_unsigned( 119,8)),
			6355 => std_logic_vector(to_unsigned( 153,8)),
			6356 => std_logic_vector(to_unsigned( 168,8)),
			6357 => std_logic_vector(to_unsigned( 192,8)),
			6358 => std_logic_vector(to_unsigned( 147,8)),
			6359 => std_logic_vector(to_unsigned( 104,8)),
			6360 => std_logic_vector(to_unsigned( 108,8)),
			6361 => std_logic_vector(to_unsigned( 214,8)),
			6362 => std_logic_vector(to_unsigned( 73,8)),
			6363 => std_logic_vector(to_unsigned( 63,8)),
			6364 => std_logic_vector(to_unsigned( 158,8)),
			6365 => std_logic_vector(to_unsigned( 187,8)),
			6366 => std_logic_vector(to_unsigned( 89,8)),
			6367 => std_logic_vector(to_unsigned( 125,8)),
			6368 => std_logic_vector(to_unsigned( 206,8)),
			6369 => std_logic_vector(to_unsigned( 92,8)),
			6370 => std_logic_vector(to_unsigned( 248,8)),
			6371 => std_logic_vector(to_unsigned( 17,8)),
			6372 => std_logic_vector(to_unsigned( 170,8)),
			6373 => std_logic_vector(to_unsigned( 59,8)),
			6374 => std_logic_vector(to_unsigned( 32,8)),
			6375 => std_logic_vector(to_unsigned( 109,8)),
			6376 => std_logic_vector(to_unsigned( 5,8)),
			6377 => std_logic_vector(to_unsigned( 0,8)),
			6378 => std_logic_vector(to_unsigned( 32,8)),
			6379 => std_logic_vector(to_unsigned( 70,8)),
			6380 => std_logic_vector(to_unsigned( 242,8)),
			6381 => std_logic_vector(to_unsigned( 176,8)),
			6382 => std_logic_vector(to_unsigned( 70,8)),
			6383 => std_logic_vector(to_unsigned( 146,8)),
			6384 => std_logic_vector(to_unsigned( 55,8)),
			6385 => std_logic_vector(to_unsigned( 56,8)),
			6386 => std_logic_vector(to_unsigned( 4,8)),
			6387 => std_logic_vector(to_unsigned( 96,8)),
			6388 => std_logic_vector(to_unsigned( 157,8)),
			6389 => std_logic_vector(to_unsigned( 203,8)),
			6390 => std_logic_vector(to_unsigned( 87,8)),
			6391 => std_logic_vector(to_unsigned( 166,8)),
			6392 => std_logic_vector(to_unsigned( 6,8)),
			6393 => std_logic_vector(to_unsigned( 51,8)),
			6394 => std_logic_vector(to_unsigned( 99,8)),
			6395 => std_logic_vector(to_unsigned( 234,8)),
			6396 => std_logic_vector(to_unsigned( 198,8)),
			6397 => std_logic_vector(to_unsigned( 42,8)),
			6398 => std_logic_vector(to_unsigned( 38,8)),
			6399 => std_logic_vector(to_unsigned( 136,8)),
			6400 => std_logic_vector(to_unsigned( 20,8)),
			6401 => std_logic_vector(to_unsigned( 156,8)),
			6402 => std_logic_vector(to_unsigned( 193,8)),
			6403 => std_logic_vector(to_unsigned( 124,8)),
			6404 => std_logic_vector(to_unsigned( 137,8)),
			6405 => std_logic_vector(to_unsigned( 225,8)),
			6406 => std_logic_vector(to_unsigned( 239,8)),
			6407 => std_logic_vector(to_unsigned( 237,8)),
			6408 => std_logic_vector(to_unsigned( 119,8)),
			6409 => std_logic_vector(to_unsigned( 254,8)),
			6410 => std_logic_vector(to_unsigned( 221,8)),
			6411 => std_logic_vector(to_unsigned( 9,8)),
			6412 => std_logic_vector(to_unsigned( 74,8)),
			6413 => std_logic_vector(to_unsigned( 218,8)),
			6414 => std_logic_vector(to_unsigned( 65,8)),
			6415 => std_logic_vector(to_unsigned( 76,8)),
			6416 => std_logic_vector(to_unsigned( 60,8)),
			6417 => std_logic_vector(to_unsigned( 86,8)),
			6418 => std_logic_vector(to_unsigned( 128,8)),
			6419 => std_logic_vector(to_unsigned( 111,8)),
			6420 => std_logic_vector(to_unsigned( 189,8)),
			6421 => std_logic_vector(to_unsigned( 246,8)),
			6422 => std_logic_vector(to_unsigned( 10,8)),
			6423 => std_logic_vector(to_unsigned( 221,8)),
			6424 => std_logic_vector(to_unsigned( 38,8)),
			6425 => std_logic_vector(to_unsigned( 254,8)),
			6426 => std_logic_vector(to_unsigned( 108,8)),
			6427 => std_logic_vector(to_unsigned( 166,8)),
			6428 => std_logic_vector(to_unsigned( 194,8)),
			6429 => std_logic_vector(to_unsigned( 144,8)),
			6430 => std_logic_vector(to_unsigned( 40,8)),
			6431 => std_logic_vector(to_unsigned( 147,8)),
			6432 => std_logic_vector(to_unsigned( 206,8)),
			6433 => std_logic_vector(to_unsigned( 50,8)),
			6434 => std_logic_vector(to_unsigned( 96,8)),
			6435 => std_logic_vector(to_unsigned( 13,8)),
			6436 => std_logic_vector(to_unsigned( 148,8)),
			6437 => std_logic_vector(to_unsigned( 214,8)),
			6438 => std_logic_vector(to_unsigned( 27,8)),
			6439 => std_logic_vector(to_unsigned( 247,8)),
			6440 => std_logic_vector(to_unsigned( 72,8)),
			6441 => std_logic_vector(to_unsigned( 83,8)),
			6442 => std_logic_vector(to_unsigned( 162,8)),
			6443 => std_logic_vector(to_unsigned( 252,8)),
			6444 => std_logic_vector(to_unsigned( 53,8)),
			6445 => std_logic_vector(to_unsigned( 66,8)),
			6446 => std_logic_vector(to_unsigned( 232,8)),
			6447 => std_logic_vector(to_unsigned( 95,8)),
			6448 => std_logic_vector(to_unsigned( 132,8)),
			6449 => std_logic_vector(to_unsigned( 224,8)),
			6450 => std_logic_vector(to_unsigned( 210,8)),
			6451 => std_logic_vector(to_unsigned( 254,8)),
			6452 => std_logic_vector(to_unsigned( 26,8)),
			6453 => std_logic_vector(to_unsigned( 127,8)),
			6454 => std_logic_vector(to_unsigned( 122,8)),
			6455 => std_logic_vector(to_unsigned( 242,8)),
			6456 => std_logic_vector(to_unsigned( 72,8)),
			6457 => std_logic_vector(to_unsigned( 237,8)),
			6458 => std_logic_vector(to_unsigned( 105,8)),
			6459 => std_logic_vector(to_unsigned( 89,8)),
			6460 => std_logic_vector(to_unsigned( 89,8)),
			6461 => std_logic_vector(to_unsigned( 147,8)),
			6462 => std_logic_vector(to_unsigned( 201,8)),
			6463 => std_logic_vector(to_unsigned( 237,8)),
			6464 => std_logic_vector(to_unsigned( 237,8)),
			6465 => std_logic_vector(to_unsigned( 50,8)),
			6466 => std_logic_vector(to_unsigned( 20,8)),
			6467 => std_logic_vector(to_unsigned( 234,8)),
			6468 => std_logic_vector(to_unsigned( 171,8)),
			6469 => std_logic_vector(to_unsigned( 51,8)),
			6470 => std_logic_vector(to_unsigned( 41,8)),
			6471 => std_logic_vector(to_unsigned( 117,8)),
			6472 => std_logic_vector(to_unsigned( 223,8)),
			6473 => std_logic_vector(to_unsigned( 89,8)),
			6474 => std_logic_vector(to_unsigned( 253,8)),
			6475 => std_logic_vector(to_unsigned( 193,8)),
			6476 => std_logic_vector(to_unsigned( 147,8)),
			6477 => std_logic_vector(to_unsigned( 155,8)),
			6478 => std_logic_vector(to_unsigned( 108,8)),
			6479 => std_logic_vector(to_unsigned( 245,8)),
			6480 => std_logic_vector(to_unsigned( 9,8)),
			6481 => std_logic_vector(to_unsigned( 64,8)),
			6482 => std_logic_vector(to_unsigned( 202,8)),
			6483 => std_logic_vector(to_unsigned( 86,8)),
			6484 => std_logic_vector(to_unsigned( 11,8)),
			6485 => std_logic_vector(to_unsigned( 210,8)),
			6486 => std_logic_vector(to_unsigned( 7,8)),
			6487 => std_logic_vector(to_unsigned( 204,8)),
			6488 => std_logic_vector(to_unsigned( 140,8)),
			6489 => std_logic_vector(to_unsigned( 77,8)),
			6490 => std_logic_vector(to_unsigned( 154,8)),
			6491 => std_logic_vector(to_unsigned( 85,8)),
			6492 => std_logic_vector(to_unsigned( 160,8)),
			6493 => std_logic_vector(to_unsigned( 71,8)),
			6494 => std_logic_vector(to_unsigned( 180,8)),
			6495 => std_logic_vector(to_unsigned( 28,8)),
			6496 => std_logic_vector(to_unsigned( 246,8)),
			6497 => std_logic_vector(to_unsigned( 32,8)),
			6498 => std_logic_vector(to_unsigned( 57,8)),
			6499 => std_logic_vector(to_unsigned( 144,8)),
			6500 => std_logic_vector(to_unsigned( 3,8)),
			6501 => std_logic_vector(to_unsigned( 36,8)),
			6502 => std_logic_vector(to_unsigned( 76,8)),
			6503 => std_logic_vector(to_unsigned( 42,8)),
			6504 => std_logic_vector(to_unsigned( 92,8)),
			6505 => std_logic_vector(to_unsigned( 191,8)),
			6506 => std_logic_vector(to_unsigned( 9,8)),
			6507 => std_logic_vector(to_unsigned( 151,8)),
			6508 => std_logic_vector(to_unsigned( 116,8)),
			6509 => std_logic_vector(to_unsigned( 121,8)),
			6510 => std_logic_vector(to_unsigned( 90,8)),
			6511 => std_logic_vector(to_unsigned( 176,8)),
			6512 => std_logic_vector(to_unsigned( 61,8)),
			6513 => std_logic_vector(to_unsigned( 18,8)),
			6514 => std_logic_vector(to_unsigned( 31,8)),
			6515 => std_logic_vector(to_unsigned( 25,8)),
			6516 => std_logic_vector(to_unsigned( 230,8)),
			6517 => std_logic_vector(to_unsigned( 164,8)),
			6518 => std_logic_vector(to_unsigned( 220,8)),
			6519 => std_logic_vector(to_unsigned( 157,8)),
			6520 => std_logic_vector(to_unsigned( 138,8)),
			6521 => std_logic_vector(to_unsigned( 227,8)),
			6522 => std_logic_vector(to_unsigned( 90,8)),
			6523 => std_logic_vector(to_unsigned( 9,8)),
			6524 => std_logic_vector(to_unsigned( 94,8)),
			6525 => std_logic_vector(to_unsigned( 59,8)),
			6526 => std_logic_vector(to_unsigned( 7,8)),
			6527 => std_logic_vector(to_unsigned( 137,8)),
			6528 => std_logic_vector(to_unsigned( 184,8)),
			6529 => std_logic_vector(to_unsigned( 211,8)),
			6530 => std_logic_vector(to_unsigned( 143,8)),
			6531 => std_logic_vector(to_unsigned( 104,8)),
			6532 => std_logic_vector(to_unsigned( 216,8)),
			6533 => std_logic_vector(to_unsigned( 55,8)),
			6534 => std_logic_vector(to_unsigned( 238,8)),
			6535 => std_logic_vector(to_unsigned( 239,8)),
			6536 => std_logic_vector(to_unsigned( 211,8)),
			6537 => std_logic_vector(to_unsigned( 171,8)),
			6538 => std_logic_vector(to_unsigned( 130,8)),
			6539 => std_logic_vector(to_unsigned( 161,8)),
			6540 => std_logic_vector(to_unsigned( 192,8)),
			6541 => std_logic_vector(to_unsigned( 143,8)),
			6542 => std_logic_vector(to_unsigned( 93,8)),
			6543 => std_logic_vector(to_unsigned( 146,8)),
			6544 => std_logic_vector(to_unsigned( 133,8)),
			6545 => std_logic_vector(to_unsigned( 17,8)),
			6546 => std_logic_vector(to_unsigned( 169,8)),
			6547 => std_logic_vector(to_unsigned( 99,8)),
			6548 => std_logic_vector(to_unsigned( 79,8)),
			6549 => std_logic_vector(to_unsigned( 160,8)),
			6550 => std_logic_vector(to_unsigned( 63,8)),
			6551 => std_logic_vector(to_unsigned( 31,8)),
			6552 => std_logic_vector(to_unsigned( 121,8)),
			6553 => std_logic_vector(to_unsigned( 106,8)),
			6554 => std_logic_vector(to_unsigned( 114,8)),
			6555 => std_logic_vector(to_unsigned( 113,8)),
			6556 => std_logic_vector(to_unsigned( 89,8)),
			6557 => std_logic_vector(to_unsigned( 48,8)),
			6558 => std_logic_vector(to_unsigned( 107,8)),
			6559 => std_logic_vector(to_unsigned( 91,8)),
			6560 => std_logic_vector(to_unsigned( 42,8)),
			6561 => std_logic_vector(to_unsigned( 31,8)),
			6562 => std_logic_vector(to_unsigned( 48,8)),
			6563 => std_logic_vector(to_unsigned( 198,8)),
			6564 => std_logic_vector(to_unsigned( 6,8)),
			6565 => std_logic_vector(to_unsigned( 225,8)),
			6566 => std_logic_vector(to_unsigned( 130,8)),
			6567 => std_logic_vector(to_unsigned( 187,8)),
			6568 => std_logic_vector(to_unsigned( 213,8)),
			6569 => std_logic_vector(to_unsigned( 173,8)),
			6570 => std_logic_vector(to_unsigned( 86,8)),
			6571 => std_logic_vector(to_unsigned( 199,8)),
			6572 => std_logic_vector(to_unsigned( 163,8)),
			6573 => std_logic_vector(to_unsigned( 90,8)),
			6574 => std_logic_vector(to_unsigned( 59,8)),
			6575 => std_logic_vector(to_unsigned( 3,8)),
			6576 => std_logic_vector(to_unsigned( 60,8)),
			6577 => std_logic_vector(to_unsigned( 114,8)),
			6578 => std_logic_vector(to_unsigned( 62,8)),
			6579 => std_logic_vector(to_unsigned( 19,8)),
			6580 => std_logic_vector(to_unsigned( 218,8)),
			6581 => std_logic_vector(to_unsigned( 233,8)),
			6582 => std_logic_vector(to_unsigned( 173,8)),
			6583 => std_logic_vector(to_unsigned( 113,8)),
			6584 => std_logic_vector(to_unsigned( 115,8)),
			6585 => std_logic_vector(to_unsigned( 148,8)),
			6586 => std_logic_vector(to_unsigned( 42,8)),
			6587 => std_logic_vector(to_unsigned( 160,8)),
			6588 => std_logic_vector(to_unsigned( 201,8)),
			6589 => std_logic_vector(to_unsigned( 110,8)),
			6590 => std_logic_vector(to_unsigned( 40,8)),
			6591 => std_logic_vector(to_unsigned( 193,8)),
			6592 => std_logic_vector(to_unsigned( 107,8)),
			6593 => std_logic_vector(to_unsigned( 102,8)),
			6594 => std_logic_vector(to_unsigned( 255,8)),
			6595 => std_logic_vector(to_unsigned( 20,8)),
			6596 => std_logic_vector(to_unsigned( 40,8)),
			6597 => std_logic_vector(to_unsigned( 204,8)),
			6598 => std_logic_vector(to_unsigned( 235,8)),
			6599 => std_logic_vector(to_unsigned( 14,8)),
			6600 => std_logic_vector(to_unsigned( 49,8)),
			6601 => std_logic_vector(to_unsigned( 234,8)),
			6602 => std_logic_vector(to_unsigned( 176,8)),
			6603 => std_logic_vector(to_unsigned( 187,8)),
			6604 => std_logic_vector(to_unsigned( 0,8)),
			6605 => std_logic_vector(to_unsigned( 162,8)),
			6606 => std_logic_vector(to_unsigned( 173,8)),
			6607 => std_logic_vector(to_unsigned( 197,8)),
			6608 => std_logic_vector(to_unsigned( 6,8)),
			6609 => std_logic_vector(to_unsigned( 228,8)),
			6610 => std_logic_vector(to_unsigned( 132,8)),
			6611 => std_logic_vector(to_unsigned( 192,8)),
			6612 => std_logic_vector(to_unsigned( 166,8)),
			6613 => std_logic_vector(to_unsigned( 228,8)),
			6614 => std_logic_vector(to_unsigned( 211,8)),
			6615 => std_logic_vector(to_unsigned( 39,8)),
			6616 => std_logic_vector(to_unsigned( 121,8)),
			6617 => std_logic_vector(to_unsigned( 153,8)),
			6618 => std_logic_vector(to_unsigned( 117,8)),
			6619 => std_logic_vector(to_unsigned( 191,8)),
			6620 => std_logic_vector(to_unsigned( 179,8)),
			6621 => std_logic_vector(to_unsigned( 23,8)),
			6622 => std_logic_vector(to_unsigned( 28,8)),
			6623 => std_logic_vector(to_unsigned( 57,8)),
			6624 => std_logic_vector(to_unsigned( 182,8)),
			6625 => std_logic_vector(to_unsigned( 234,8)),
			6626 => std_logic_vector(to_unsigned( 121,8)),
			6627 => std_logic_vector(to_unsigned( 60,8)),
			6628 => std_logic_vector(to_unsigned( 232,8)),
			6629 => std_logic_vector(to_unsigned( 15,8)),
			6630 => std_logic_vector(to_unsigned( 9,8)),
			6631 => std_logic_vector(to_unsigned( 241,8)),
			6632 => std_logic_vector(to_unsigned( 78,8)),
			6633 => std_logic_vector(to_unsigned( 134,8)),
			6634 => std_logic_vector(to_unsigned( 221,8)),
			6635 => std_logic_vector(to_unsigned( 29,8)),
			6636 => std_logic_vector(to_unsigned( 144,8)),
			6637 => std_logic_vector(to_unsigned( 109,8)),
			6638 => std_logic_vector(to_unsigned( 51,8)),
			6639 => std_logic_vector(to_unsigned( 71,8)),
			6640 => std_logic_vector(to_unsigned( 248,8)),
			6641 => std_logic_vector(to_unsigned( 11,8)),
			6642 => std_logic_vector(to_unsigned( 171,8)),
			6643 => std_logic_vector(to_unsigned( 84,8)),
			6644 => std_logic_vector(to_unsigned( 162,8)),
			6645 => std_logic_vector(to_unsigned( 231,8)),
			6646 => std_logic_vector(to_unsigned( 30,8)),
			6647 => std_logic_vector(to_unsigned( 214,8)),
			6648 => std_logic_vector(to_unsigned( 196,8)),
			6649 => std_logic_vector(to_unsigned( 116,8)),
			6650 => std_logic_vector(to_unsigned( 230,8)),
			6651 => std_logic_vector(to_unsigned( 179,8)),
			6652 => std_logic_vector(to_unsigned( 22,8)),
			6653 => std_logic_vector(to_unsigned( 229,8)),
			6654 => std_logic_vector(to_unsigned( 238,8)),
			6655 => std_logic_vector(to_unsigned( 133,8)),
			6656 => std_logic_vector(to_unsigned( 115,8)),
			6657 => std_logic_vector(to_unsigned( 254,8)),
			6658 => std_logic_vector(to_unsigned( 241,8)),
			6659 => std_logic_vector(to_unsigned( 178,8)),
			6660 => std_logic_vector(to_unsigned( 139,8)),
			6661 => std_logic_vector(to_unsigned( 78,8)),
			6662 => std_logic_vector(to_unsigned( 214,8)),
			6663 => std_logic_vector(to_unsigned( 21,8)),
			6664 => std_logic_vector(to_unsigned( 174,8)),
			6665 => std_logic_vector(to_unsigned( 139,8)),
			6666 => std_logic_vector(to_unsigned( 152,8)),
			6667 => std_logic_vector(to_unsigned( 250,8)),
			6668 => std_logic_vector(to_unsigned( 229,8)),
			6669 => std_logic_vector(to_unsigned( 39,8)),
			6670 => std_logic_vector(to_unsigned( 138,8)),
			6671 => std_logic_vector(to_unsigned( 203,8)),
			6672 => std_logic_vector(to_unsigned( 222,8)),
			6673 => std_logic_vector(to_unsigned( 193,8)),
			6674 => std_logic_vector(to_unsigned( 206,8)),
			6675 => std_logic_vector(to_unsigned( 67,8)),
			6676 => std_logic_vector(to_unsigned( 245,8)),
			6677 => std_logic_vector(to_unsigned( 161,8)),
			6678 => std_logic_vector(to_unsigned( 31,8)),
			6679 => std_logic_vector(to_unsigned( 87,8)),
			6680 => std_logic_vector(to_unsigned( 166,8)),
			6681 => std_logic_vector(to_unsigned( 150,8)),
			6682 => std_logic_vector(to_unsigned( 162,8)),
			6683 => std_logic_vector(to_unsigned( 36,8)),
			6684 => std_logic_vector(to_unsigned( 83,8)),
			6685 => std_logic_vector(to_unsigned( 102,8)),
			6686 => std_logic_vector(to_unsigned( 56,8)),
			6687 => std_logic_vector(to_unsigned( 140,8)),
			6688 => std_logic_vector(to_unsigned( 253,8)),
			6689 => std_logic_vector(to_unsigned( 138,8)),
			6690 => std_logic_vector(to_unsigned( 195,8)),
			6691 => std_logic_vector(to_unsigned( 40,8)),
			6692 => std_logic_vector(to_unsigned( 126,8)),
			6693 => std_logic_vector(to_unsigned( 106,8)),
			6694 => std_logic_vector(to_unsigned( 198,8)),
			6695 => std_logic_vector(to_unsigned( 54,8)),
			6696 => std_logic_vector(to_unsigned( 183,8)),
			6697 => std_logic_vector(to_unsigned( 73,8)),
			6698 => std_logic_vector(to_unsigned( 120,8)),
			6699 => std_logic_vector(to_unsigned( 222,8)),
			6700 => std_logic_vector(to_unsigned( 112,8)),
			6701 => std_logic_vector(to_unsigned( 107,8)),
			6702 => std_logic_vector(to_unsigned( 160,8)),
			6703 => std_logic_vector(to_unsigned( 17,8)),
			6704 => std_logic_vector(to_unsigned( 186,8)),
			6705 => std_logic_vector(to_unsigned( 54,8)),
			6706 => std_logic_vector(to_unsigned( 71,8)),
			6707 => std_logic_vector(to_unsigned( 180,8)),
			6708 => std_logic_vector(to_unsigned( 5,8)),
			6709 => std_logic_vector(to_unsigned( 44,8)),
			6710 => std_logic_vector(to_unsigned( 16,8)),
			6711 => std_logic_vector(to_unsigned( 67,8)),
			6712 => std_logic_vector(to_unsigned( 169,8)),
			6713 => std_logic_vector(to_unsigned( 146,8)),
			6714 => std_logic_vector(to_unsigned( 68,8)),
			6715 => std_logic_vector(to_unsigned( 12,8)),
			6716 => std_logic_vector(to_unsigned( 221,8)),
			6717 => std_logic_vector(to_unsigned( 60,8)),
			6718 => std_logic_vector(to_unsigned( 161,8)),
			6719 => std_logic_vector(to_unsigned( 219,8)),
			6720 => std_logic_vector(to_unsigned( 97,8)),
			6721 => std_logic_vector(to_unsigned( 219,8)),
			6722 => std_logic_vector(to_unsigned( 19,8)),
			6723 => std_logic_vector(to_unsigned( 161,8)),
			6724 => std_logic_vector(to_unsigned( 162,8)),
			6725 => std_logic_vector(to_unsigned( 117,8)),
			6726 => std_logic_vector(to_unsigned( 170,8)),
			6727 => std_logic_vector(to_unsigned( 146,8)),
			6728 => std_logic_vector(to_unsigned( 128,8)),
			6729 => std_logic_vector(to_unsigned( 34,8)),
			6730 => std_logic_vector(to_unsigned( 197,8)),
			6731 => std_logic_vector(to_unsigned( 70,8)),
			6732 => std_logic_vector(to_unsigned( 84,8)),
			6733 => std_logic_vector(to_unsigned( 84,8)),
			6734 => std_logic_vector(to_unsigned( 189,8)),
			6735 => std_logic_vector(to_unsigned( 25,8)),
			6736 => std_logic_vector(to_unsigned( 194,8)),
			6737 => std_logic_vector(to_unsigned( 143,8)),
			6738 => std_logic_vector(to_unsigned( 49,8)),
			6739 => std_logic_vector(to_unsigned( 144,8)),
			6740 => std_logic_vector(to_unsigned( 178,8)),
			6741 => std_logic_vector(to_unsigned( 185,8)),
			6742 => std_logic_vector(to_unsigned( 229,8)),
			6743 => std_logic_vector(to_unsigned( 30,8)),
			6744 => std_logic_vector(to_unsigned( 111,8)),
			6745 => std_logic_vector(to_unsigned( 218,8)),
			6746 => std_logic_vector(to_unsigned( 175,8)),
			6747 => std_logic_vector(to_unsigned( 19,8)),
			6748 => std_logic_vector(to_unsigned( 115,8)),
			6749 => std_logic_vector(to_unsigned( 253,8)),
			6750 => std_logic_vector(to_unsigned( 227,8)),
			6751 => std_logic_vector(to_unsigned( 226,8)),
			6752 => std_logic_vector(to_unsigned( 217,8)),
			6753 => std_logic_vector(to_unsigned( 75,8)),
			6754 => std_logic_vector(to_unsigned( 38,8)),
			6755 => std_logic_vector(to_unsigned( 133,8)),
			6756 => std_logic_vector(to_unsigned( 93,8)),
			6757 => std_logic_vector(to_unsigned( 201,8)),
			6758 => std_logic_vector(to_unsigned( 241,8)),
			6759 => std_logic_vector(to_unsigned( 66,8)),
			6760 => std_logic_vector(to_unsigned( 208,8)),
			6761 => std_logic_vector(to_unsigned( 224,8)),
			6762 => std_logic_vector(to_unsigned( 123,8)),
			6763 => std_logic_vector(to_unsigned( 65,8)),
			6764 => std_logic_vector(to_unsigned( 90,8)),
			6765 => std_logic_vector(to_unsigned( 78,8)),
			6766 => std_logic_vector(to_unsigned( 146,8)),
			6767 => std_logic_vector(to_unsigned( 170,8)),
			6768 => std_logic_vector(to_unsigned( 226,8)),
			6769 => std_logic_vector(to_unsigned( 176,8)),
			6770 => std_logic_vector(to_unsigned( 221,8)),
			6771 => std_logic_vector(to_unsigned( 113,8)),
			6772 => std_logic_vector(to_unsigned( 28,8)),
			6773 => std_logic_vector(to_unsigned( 193,8)),
			6774 => std_logic_vector(to_unsigned( 157,8)),
			6775 => std_logic_vector(to_unsigned( 78,8)),
			6776 => std_logic_vector(to_unsigned( 28,8)),
			6777 => std_logic_vector(to_unsigned( 211,8)),
			6778 => std_logic_vector(to_unsigned( 43,8)),
			6779 => std_logic_vector(to_unsigned( 172,8)),
			6780 => std_logic_vector(to_unsigned( 94,8)),
			6781 => std_logic_vector(to_unsigned( 29,8)),
			6782 => std_logic_vector(to_unsigned( 110,8)),
			6783 => std_logic_vector(to_unsigned( 57,8)),
			6784 => std_logic_vector(to_unsigned( 38,8)),
			6785 => std_logic_vector(to_unsigned( 109,8)),
			6786 => std_logic_vector(to_unsigned( 139,8)),
			6787 => std_logic_vector(to_unsigned( 242,8)),
			6788 => std_logic_vector(to_unsigned( 235,8)),
			6789 => std_logic_vector(to_unsigned( 36,8)),
			6790 => std_logic_vector(to_unsigned( 90,8)),
			6791 => std_logic_vector(to_unsigned( 156,8)),
			6792 => std_logic_vector(to_unsigned( 74,8)),
			6793 => std_logic_vector(to_unsigned( 31,8)),
			6794 => std_logic_vector(to_unsigned( 117,8)),
			6795 => std_logic_vector(to_unsigned( 73,8)),
			6796 => std_logic_vector(to_unsigned( 109,8)),
			6797 => std_logic_vector(to_unsigned( 180,8)),
			6798 => std_logic_vector(to_unsigned( 120,8)),
			6799 => std_logic_vector(to_unsigned( 187,8)),
			6800 => std_logic_vector(to_unsigned( 42,8)),
			6801 => std_logic_vector(to_unsigned( 149,8)),
			6802 => std_logic_vector(to_unsigned( 183,8)),
			6803 => std_logic_vector(to_unsigned( 135,8)),
			6804 => std_logic_vector(to_unsigned( 17,8)),
			6805 => std_logic_vector(to_unsigned( 86,8)),
			6806 => std_logic_vector(to_unsigned( 7,8)),
			6807 => std_logic_vector(to_unsigned( 217,8)),
			6808 => std_logic_vector(to_unsigned( 124,8)),
			6809 => std_logic_vector(to_unsigned( 70,8)),
			6810 => std_logic_vector(to_unsigned( 24,8)),
			6811 => std_logic_vector(to_unsigned( 35,8)),
			6812 => std_logic_vector(to_unsigned( 139,8)),
			6813 => std_logic_vector(to_unsigned( 240,8)),
			6814 => std_logic_vector(to_unsigned( 53,8)),
			6815 => std_logic_vector(to_unsigned( 86,8)),
			6816 => std_logic_vector(to_unsigned( 174,8)),
			6817 => std_logic_vector(to_unsigned( 255,8)),
			6818 => std_logic_vector(to_unsigned( 106,8)),
			6819 => std_logic_vector(to_unsigned( 143,8)),
			6820 => std_logic_vector(to_unsigned( 24,8)),
			6821 => std_logic_vector(to_unsigned( 216,8)),
			6822 => std_logic_vector(to_unsigned( 56,8)),
			6823 => std_logic_vector(to_unsigned( 118,8)),
			6824 => std_logic_vector(to_unsigned( 136,8)),
			6825 => std_logic_vector(to_unsigned( 182,8)),
			6826 => std_logic_vector(to_unsigned( 43,8)),
			6827 => std_logic_vector(to_unsigned( 127,8)),
			6828 => std_logic_vector(to_unsigned( 201,8)),
			6829 => std_logic_vector(to_unsigned( 199,8)),
			6830 => std_logic_vector(to_unsigned( 90,8)),
			6831 => std_logic_vector(to_unsigned( 172,8)),
			6832 => std_logic_vector(to_unsigned( 198,8)),
			6833 => std_logic_vector(to_unsigned( 25,8)),
			6834 => std_logic_vector(to_unsigned( 72,8)),
			6835 => std_logic_vector(to_unsigned( 79,8)),
			6836 => std_logic_vector(to_unsigned( 27,8)),
			6837 => std_logic_vector(to_unsigned( 240,8)),
			6838 => std_logic_vector(to_unsigned( 192,8)),
			6839 => std_logic_vector(to_unsigned( 107,8)),
			6840 => std_logic_vector(to_unsigned( 145,8)),
			6841 => std_logic_vector(to_unsigned( 21,8)),
			6842 => std_logic_vector(to_unsigned( 202,8)),
			6843 => std_logic_vector(to_unsigned( 40,8)),
			6844 => std_logic_vector(to_unsigned( 125,8)),
			6845 => std_logic_vector(to_unsigned( 181,8)),
			6846 => std_logic_vector(to_unsigned( 61,8)),
			6847 => std_logic_vector(to_unsigned( 202,8)),
			6848 => std_logic_vector(to_unsigned( 14,8)),
			6849 => std_logic_vector(to_unsigned( 37,8)),
			6850 => std_logic_vector(to_unsigned( 133,8)),
			6851 => std_logic_vector(to_unsigned( 229,8)),
			6852 => std_logic_vector(to_unsigned( 0,8)),
			6853 => std_logic_vector(to_unsigned( 225,8)),
			6854 => std_logic_vector(to_unsigned( 184,8)),
			6855 => std_logic_vector(to_unsigned( 142,8)),
			6856 => std_logic_vector(to_unsigned( 106,8)),
			6857 => std_logic_vector(to_unsigned( 214,8)),
			6858 => std_logic_vector(to_unsigned( 64,8)),
			6859 => std_logic_vector(to_unsigned( 6,8)),
			6860 => std_logic_vector(to_unsigned( 111,8)),
			6861 => std_logic_vector(to_unsigned( 217,8)),
			6862 => std_logic_vector(to_unsigned( 211,8)),
			6863 => std_logic_vector(to_unsigned( 2,8)),
			6864 => std_logic_vector(to_unsigned( 120,8)),
			6865 => std_logic_vector(to_unsigned( 216,8)),
			6866 => std_logic_vector(to_unsigned( 24,8)),
			6867 => std_logic_vector(to_unsigned( 39,8)),
			6868 => std_logic_vector(to_unsigned( 157,8)),
			6869 => std_logic_vector(to_unsigned( 127,8)),
			6870 => std_logic_vector(to_unsigned( 129,8)),
			6871 => std_logic_vector(to_unsigned( 199,8)),
			6872 => std_logic_vector(to_unsigned( 80,8)),
			6873 => std_logic_vector(to_unsigned( 163,8)),
			6874 => std_logic_vector(to_unsigned( 2,8)),
			6875 => std_logic_vector(to_unsigned( 207,8)),
			6876 => std_logic_vector(to_unsigned( 158,8)),
			6877 => std_logic_vector(to_unsigned( 117,8)),
			6878 => std_logic_vector(to_unsigned( 155,8)),
			6879 => std_logic_vector(to_unsigned( 231,8)),
			6880 => std_logic_vector(to_unsigned( 164,8)),
			6881 => std_logic_vector(to_unsigned( 99,8)),
			6882 => std_logic_vector(to_unsigned( 139,8)),
			6883 => std_logic_vector(to_unsigned( 4,8)),
			6884 => std_logic_vector(to_unsigned( 187,8)),
			6885 => std_logic_vector(to_unsigned( 49,8)),
			6886 => std_logic_vector(to_unsigned( 184,8)),
			6887 => std_logic_vector(to_unsigned( 242,8)),
			6888 => std_logic_vector(to_unsigned( 237,8)),
			6889 => std_logic_vector(to_unsigned( 39,8)),
			6890 => std_logic_vector(to_unsigned( 205,8)),
			6891 => std_logic_vector(to_unsigned( 112,8)),
			6892 => std_logic_vector(to_unsigned( 22,8)),
			6893 => std_logic_vector(to_unsigned( 206,8)),
			6894 => std_logic_vector(to_unsigned( 184,8)),
			6895 => std_logic_vector(to_unsigned( 119,8)),
			6896 => std_logic_vector(to_unsigned( 49,8)),
			6897 => std_logic_vector(to_unsigned( 88,8)),
			6898 => std_logic_vector(to_unsigned( 136,8)),
			6899 => std_logic_vector(to_unsigned( 16,8)),
			6900 => std_logic_vector(to_unsigned( 171,8)),
			6901 => std_logic_vector(to_unsigned( 164,8)),
			6902 => std_logic_vector(to_unsigned( 145,8)),
			6903 => std_logic_vector(to_unsigned( 206,8)),
			6904 => std_logic_vector(to_unsigned( 131,8)),
			6905 => std_logic_vector(to_unsigned( 33,8)),
			6906 => std_logic_vector(to_unsigned( 169,8)),
			6907 => std_logic_vector(to_unsigned( 220,8)),
			6908 => std_logic_vector(to_unsigned( 149,8)),
			6909 => std_logic_vector(to_unsigned( 162,8)),
			6910 => std_logic_vector(to_unsigned( 237,8)),
			6911 => std_logic_vector(to_unsigned( 240,8)),
			6912 => std_logic_vector(to_unsigned( 188,8)),
			6913 => std_logic_vector(to_unsigned( 96,8)),
			6914 => std_logic_vector(to_unsigned( 136,8)),
			6915 => std_logic_vector(to_unsigned( 111,8)),
			6916 => std_logic_vector(to_unsigned( 177,8)),
			6917 => std_logic_vector(to_unsigned( 160,8)),
			6918 => std_logic_vector(to_unsigned( 167,8)),
			6919 => std_logic_vector(to_unsigned( 245,8)),
			6920 => std_logic_vector(to_unsigned( 95,8)),
			6921 => std_logic_vector(to_unsigned( 202,8)),
			6922 => std_logic_vector(to_unsigned( 94,8)),
			6923 => std_logic_vector(to_unsigned( 36,8)),
			6924 => std_logic_vector(to_unsigned( 8,8)),
			6925 => std_logic_vector(to_unsigned( 143,8)),
			6926 => std_logic_vector(to_unsigned( 165,8)),
			6927 => std_logic_vector(to_unsigned( 88,8)),
			6928 => std_logic_vector(to_unsigned( 54,8)),
			6929 => std_logic_vector(to_unsigned( 5,8)),
			6930 => std_logic_vector(to_unsigned( 106,8)),
			6931 => std_logic_vector(to_unsigned( 61,8)),
			6932 => std_logic_vector(to_unsigned( 71,8)),
			6933 => std_logic_vector(to_unsigned( 235,8)),
			6934 => std_logic_vector(to_unsigned( 39,8)),
			6935 => std_logic_vector(to_unsigned( 69,8)),
			6936 => std_logic_vector(to_unsigned( 101,8)),
			6937 => std_logic_vector(to_unsigned( 196,8)),
			6938 => std_logic_vector(to_unsigned( 127,8)),
			6939 => std_logic_vector(to_unsigned( 20,8)),
			6940 => std_logic_vector(to_unsigned( 104,8)),
			6941 => std_logic_vector(to_unsigned( 95,8)),
			6942 => std_logic_vector(to_unsigned( 230,8)),
			6943 => std_logic_vector(to_unsigned( 150,8)),
			6944 => std_logic_vector(to_unsigned( 186,8)),
			6945 => std_logic_vector(to_unsigned( 255,8)),
			6946 => std_logic_vector(to_unsigned( 243,8)),
			6947 => std_logic_vector(to_unsigned( 149,8)),
			6948 => std_logic_vector(to_unsigned( 219,8)),
			6949 => std_logic_vector(to_unsigned( 24,8)),
			6950 => std_logic_vector(to_unsigned( 8,8)),
			6951 => std_logic_vector(to_unsigned( 24,8)),
			6952 => std_logic_vector(to_unsigned( 67,8)),
			6953 => std_logic_vector(to_unsigned( 108,8)),
			6954 => std_logic_vector(to_unsigned( 3,8)),
			6955 => std_logic_vector(to_unsigned( 121,8)),
			6956 => std_logic_vector(to_unsigned( 189,8)),
			6957 => std_logic_vector(to_unsigned( 42,8)),
			6958 => std_logic_vector(to_unsigned( 199,8)),
			6959 => std_logic_vector(to_unsigned( 179,8)),
			6960 => std_logic_vector(to_unsigned( 126,8)),
			6961 => std_logic_vector(to_unsigned( 187,8)),
			6962 => std_logic_vector(to_unsigned( 223,8)),
			6963 => std_logic_vector(to_unsigned( 92,8)),
			6964 => std_logic_vector(to_unsigned( 174,8)),
			6965 => std_logic_vector(to_unsigned( 51,8)),
			6966 => std_logic_vector(to_unsigned( 65,8)),
			6967 => std_logic_vector(to_unsigned( 222,8)),
			6968 => std_logic_vector(to_unsigned( 234,8)),
			6969 => std_logic_vector(to_unsigned( 96,8)),
			6970 => std_logic_vector(to_unsigned( 219,8)),
			6971 => std_logic_vector(to_unsigned( 183,8)),
			6972 => std_logic_vector(to_unsigned( 249,8)),
			6973 => std_logic_vector(to_unsigned( 150,8)),
			6974 => std_logic_vector(to_unsigned( 146,8)),
			6975 => std_logic_vector(to_unsigned( 208,8)),
			6976 => std_logic_vector(to_unsigned( 5,8)),
			6977 => std_logic_vector(to_unsigned( 156,8)),
			6978 => std_logic_vector(to_unsigned( 189,8)),
			6979 => std_logic_vector(to_unsigned( 131,8)),
			6980 => std_logic_vector(to_unsigned( 182,8)),
			6981 => std_logic_vector(to_unsigned( 13,8)),
			6982 => std_logic_vector(to_unsigned( 84,8)),
			6983 => std_logic_vector(to_unsigned( 162,8)),
			6984 => std_logic_vector(to_unsigned( 240,8)),
			6985 => std_logic_vector(to_unsigned( 220,8)),
			6986 => std_logic_vector(to_unsigned( 59,8)),
			6987 => std_logic_vector(to_unsigned( 167,8)),
			6988 => std_logic_vector(to_unsigned( 82,8)),
			6989 => std_logic_vector(to_unsigned( 227,8)),
			6990 => std_logic_vector(to_unsigned( 251,8)),
			6991 => std_logic_vector(to_unsigned( 26,8)),
			6992 => std_logic_vector(to_unsigned( 28,8)),
			6993 => std_logic_vector(to_unsigned( 95,8)),
			6994 => std_logic_vector(to_unsigned( 44,8)),
			6995 => std_logic_vector(to_unsigned( 230,8)),
			6996 => std_logic_vector(to_unsigned( 7,8)),
			6997 => std_logic_vector(to_unsigned( 135,8)),
			6998 => std_logic_vector(to_unsigned( 30,8)),
			6999 => std_logic_vector(to_unsigned( 124,8)),
			7000 => std_logic_vector(to_unsigned( 12,8)),
			7001 => std_logic_vector(to_unsigned( 164,8)),
			7002 => std_logic_vector(to_unsigned( 91,8)),
			7003 => std_logic_vector(to_unsigned( 175,8)),
			7004 => std_logic_vector(to_unsigned( 187,8)),
			7005 => std_logic_vector(to_unsigned( 118,8)),
			7006 => std_logic_vector(to_unsigned( 59,8)),
			7007 => std_logic_vector(to_unsigned( 203,8)),
			7008 => std_logic_vector(to_unsigned( 172,8)),
			7009 => std_logic_vector(to_unsigned( 135,8)),
			7010 => std_logic_vector(to_unsigned( 155,8)),
			7011 => std_logic_vector(to_unsigned( 214,8)),
			7012 => std_logic_vector(to_unsigned( 146,8)),
			7013 => std_logic_vector(to_unsigned( 30,8)),
			7014 => std_logic_vector(to_unsigned( 107,8)),
			7015 => std_logic_vector(to_unsigned( 169,8)),
			7016 => std_logic_vector(to_unsigned( 156,8)),
			7017 => std_logic_vector(to_unsigned( 72,8)),
			7018 => std_logic_vector(to_unsigned( 111,8)),
			7019 => std_logic_vector(to_unsigned( 110,8)),
			7020 => std_logic_vector(to_unsigned( 157,8)),
			7021 => std_logic_vector(to_unsigned( 224,8)),
			7022 => std_logic_vector(to_unsigned( 176,8)),
			7023 => std_logic_vector(to_unsigned( 29,8)),
			7024 => std_logic_vector(to_unsigned( 60,8)),
			7025 => std_logic_vector(to_unsigned( 155,8)),
			7026 => std_logic_vector(to_unsigned( 198,8)),
			7027 => std_logic_vector(to_unsigned( 1,8)),
			7028 => std_logic_vector(to_unsigned( 15,8)),
			7029 => std_logic_vector(to_unsigned( 48,8)),
			7030 => std_logic_vector(to_unsigned( 68,8)),
			7031 => std_logic_vector(to_unsigned( 40,8)),
			7032 => std_logic_vector(to_unsigned( 63,8)),
			7033 => std_logic_vector(to_unsigned( 211,8)),
			7034 => std_logic_vector(to_unsigned( 66,8)),
			7035 => std_logic_vector(to_unsigned( 41,8)),
			7036 => std_logic_vector(to_unsigned( 114,8)),
			7037 => std_logic_vector(to_unsigned( 0,8)),
			7038 => std_logic_vector(to_unsigned( 86,8)),
			7039 => std_logic_vector(to_unsigned( 238,8)),
			7040 => std_logic_vector(to_unsigned( 208,8)),
			7041 => std_logic_vector(to_unsigned( 243,8)),
			7042 => std_logic_vector(to_unsigned( 239,8)),
			7043 => std_logic_vector(to_unsigned( 132,8)),
			7044 => std_logic_vector(to_unsigned( 250,8)),
			7045 => std_logic_vector(to_unsigned( 245,8)),
			7046 => std_logic_vector(to_unsigned( 58,8)),
			7047 => std_logic_vector(to_unsigned( 176,8)),
			7048 => std_logic_vector(to_unsigned( 38,8)),
			7049 => std_logic_vector(to_unsigned( 253,8)),
			7050 => std_logic_vector(to_unsigned( 209,8)),
			7051 => std_logic_vector(to_unsigned( 247,8)),
			7052 => std_logic_vector(to_unsigned( 46,8)),
			7053 => std_logic_vector(to_unsigned( 28,8)),
			7054 => std_logic_vector(to_unsigned( 49,8)),
			7055 => std_logic_vector(to_unsigned( 128,8)),
			7056 => std_logic_vector(to_unsigned( 241,8)),
			7057 => std_logic_vector(to_unsigned( 193,8)),
			7058 => std_logic_vector(to_unsigned( 234,8)),
			7059 => std_logic_vector(to_unsigned( 48,8)),
			7060 => std_logic_vector(to_unsigned( 158,8)),
			7061 => std_logic_vector(to_unsigned( 158,8)),
			7062 => std_logic_vector(to_unsigned( 160,8)),
			7063 => std_logic_vector(to_unsigned( 153,8)),
			7064 => std_logic_vector(to_unsigned( 100,8)),
			7065 => std_logic_vector(to_unsigned( 255,8)),
			7066 => std_logic_vector(to_unsigned( 175,8)),
			7067 => std_logic_vector(to_unsigned( 178,8)),
			7068 => std_logic_vector(to_unsigned( 140,8)),
			7069 => std_logic_vector(to_unsigned( 240,8)),
			7070 => std_logic_vector(to_unsigned( 8,8)),
			7071 => std_logic_vector(to_unsigned( 115,8)),
			7072 => std_logic_vector(to_unsigned( 3,8)),
			7073 => std_logic_vector(to_unsigned( 236,8)),
			7074 => std_logic_vector(to_unsigned( 83,8)),
			7075 => std_logic_vector(to_unsigned( 63,8)),
			7076 => std_logic_vector(to_unsigned( 42,8)),
			7077 => std_logic_vector(to_unsigned( 18,8)),
			7078 => std_logic_vector(to_unsigned( 224,8)),
			7079 => std_logic_vector(to_unsigned( 143,8)),
			7080 => std_logic_vector(to_unsigned( 160,8)),
			7081 => std_logic_vector(to_unsigned( 137,8)),
			7082 => std_logic_vector(to_unsigned( 189,8)),
			7083 => std_logic_vector(to_unsigned( 126,8)),
			7084 => std_logic_vector(to_unsigned( 7,8)),
			7085 => std_logic_vector(to_unsigned( 23,8)),
			7086 => std_logic_vector(to_unsigned( 145,8)),
			7087 => std_logic_vector(to_unsigned( 158,8)),
			7088 => std_logic_vector(to_unsigned( 222,8)),
			7089 => std_logic_vector(to_unsigned( 33,8)),
			7090 => std_logic_vector(to_unsigned( 204,8)),
			7091 => std_logic_vector(to_unsigned( 3,8)),
			7092 => std_logic_vector(to_unsigned( 207,8)),
			7093 => std_logic_vector(to_unsigned( 35,8)),
			7094 => std_logic_vector(to_unsigned( 103,8)),
			7095 => std_logic_vector(to_unsigned( 165,8)),
			7096 => std_logic_vector(to_unsigned( 45,8)),
			7097 => std_logic_vector(to_unsigned( 43,8)),
			7098 => std_logic_vector(to_unsigned( 107,8)),
			7099 => std_logic_vector(to_unsigned( 130,8)),
			7100 => std_logic_vector(to_unsigned( 96,8)),
			7101 => std_logic_vector(to_unsigned( 210,8)),
			7102 => std_logic_vector(to_unsigned( 53,8)),
			7103 => std_logic_vector(to_unsigned( 46,8)),
			7104 => std_logic_vector(to_unsigned( 139,8)),
			7105 => std_logic_vector(to_unsigned( 231,8)),
			7106 => std_logic_vector(to_unsigned( 120,8)),
			7107 => std_logic_vector(to_unsigned( 169,8)),
			7108 => std_logic_vector(to_unsigned( 112,8)),
			7109 => std_logic_vector(to_unsigned( 55,8)),
			7110 => std_logic_vector(to_unsigned( 43,8)),
			7111 => std_logic_vector(to_unsigned( 88,8)),
			7112 => std_logic_vector(to_unsigned( 119,8)),
			7113 => std_logic_vector(to_unsigned( 131,8)),
			7114 => std_logic_vector(to_unsigned( 18,8)),
			7115 => std_logic_vector(to_unsigned( 154,8)),
			7116 => std_logic_vector(to_unsigned( 109,8)),
			7117 => std_logic_vector(to_unsigned( 162,8)),
			7118 => std_logic_vector(to_unsigned( 94,8)),
			7119 => std_logic_vector(to_unsigned( 189,8)),
			7120 => std_logic_vector(to_unsigned( 71,8)),
			7121 => std_logic_vector(to_unsigned( 64,8)),
			7122 => std_logic_vector(to_unsigned( 238,8)),
			7123 => std_logic_vector(to_unsigned( 32,8)),
			7124 => std_logic_vector(to_unsigned( 89,8)),
			7125 => std_logic_vector(to_unsigned( 14,8)),
			7126 => std_logic_vector(to_unsigned( 111,8)),
			7127 => std_logic_vector(to_unsigned( 95,8)),
			7128 => std_logic_vector(to_unsigned( 163,8)),
			7129 => std_logic_vector(to_unsigned( 208,8)),
			7130 => std_logic_vector(to_unsigned( 32,8)),
			7131 => std_logic_vector(to_unsigned( 123,8)),
			7132 => std_logic_vector(to_unsigned( 69,8)),
			7133 => std_logic_vector(to_unsigned( 228,8)),
			7134 => std_logic_vector(to_unsigned( 117,8)),
			7135 => std_logic_vector(to_unsigned( 106,8)),
			7136 => std_logic_vector(to_unsigned( 237,8)),
			7137 => std_logic_vector(to_unsigned( 127,8)),
			7138 => std_logic_vector(to_unsigned( 228,8)),
			7139 => std_logic_vector(to_unsigned( 214,8)),
			7140 => std_logic_vector(to_unsigned( 80,8)),
			7141 => std_logic_vector(to_unsigned( 74,8)),
			7142 => std_logic_vector(to_unsigned( 50,8)),
			7143 => std_logic_vector(to_unsigned( 15,8)),
			7144 => std_logic_vector(to_unsigned( 27,8)),
			7145 => std_logic_vector(to_unsigned( 162,8)),
			7146 => std_logic_vector(to_unsigned( 18,8)),
			7147 => std_logic_vector(to_unsigned( 247,8)),
			7148 => std_logic_vector(to_unsigned( 104,8)),
			7149 => std_logic_vector(to_unsigned( 229,8)),
			7150 => std_logic_vector(to_unsigned( 247,8)),
			7151 => std_logic_vector(to_unsigned( 177,8)),
			7152 => std_logic_vector(to_unsigned( 179,8)),
			7153 => std_logic_vector(to_unsigned( 216,8)),
			7154 => std_logic_vector(to_unsigned( 18,8)),
			7155 => std_logic_vector(to_unsigned( 22,8)),
			7156 => std_logic_vector(to_unsigned( 154,8)),
			7157 => std_logic_vector(to_unsigned( 85,8)),
			7158 => std_logic_vector(to_unsigned( 221,8)),
			7159 => std_logic_vector(to_unsigned( 40,8)),
			7160 => std_logic_vector(to_unsigned( 161,8)),
			7161 => std_logic_vector(to_unsigned( 109,8)),
			7162 => std_logic_vector(to_unsigned( 82,8)),
			7163 => std_logic_vector(to_unsigned( 41,8)),
			7164 => std_logic_vector(to_unsigned( 69,8)),
			7165 => std_logic_vector(to_unsigned( 93,8)),
			7166 => std_logic_vector(to_unsigned( 233,8)),
			7167 => std_logic_vector(to_unsigned( 18,8)),
			7168 => std_logic_vector(to_unsigned( 184,8)),
			7169 => std_logic_vector(to_unsigned( 250,8)),
			7170 => std_logic_vector(to_unsigned( 71,8)),
			7171 => std_logic_vector(to_unsigned( 198,8)),
			7172 => std_logic_vector(to_unsigned( 188,8)),
			7173 => std_logic_vector(to_unsigned( 27,8)),
			7174 => std_logic_vector(to_unsigned( 186,8)),
			7175 => std_logic_vector(to_unsigned( 221,8)),
			7176 => std_logic_vector(to_unsigned( 36,8)),
			7177 => std_logic_vector(to_unsigned( 189,8)),
			7178 => std_logic_vector(to_unsigned( 90,8)),
			7179 => std_logic_vector(to_unsigned( 249,8)),
			7180 => std_logic_vector(to_unsigned( 249,8)),
			7181 => std_logic_vector(to_unsigned( 238,8)),
			7182 => std_logic_vector(to_unsigned( 141,8)),
			7183 => std_logic_vector(to_unsigned( 190,8)),
			7184 => std_logic_vector(to_unsigned( 210,8)),
			7185 => std_logic_vector(to_unsigned( 28,8)),
			7186 => std_logic_vector(to_unsigned( 58,8)),
			7187 => std_logic_vector(to_unsigned( 39,8)),
			7188 => std_logic_vector(to_unsigned( 56,8)),
			7189 => std_logic_vector(to_unsigned( 96,8)),
			7190 => std_logic_vector(to_unsigned( 198,8)),
			7191 => std_logic_vector(to_unsigned( 52,8)),
			7192 => std_logic_vector(to_unsigned( 31,8)),
			7193 => std_logic_vector(to_unsigned( 48,8)),
			7194 => std_logic_vector(to_unsigned( 164,8)),
			7195 => std_logic_vector(to_unsigned( 165,8)),
			7196 => std_logic_vector(to_unsigned( 210,8)),
			7197 => std_logic_vector(to_unsigned( 138,8)),
			7198 => std_logic_vector(to_unsigned( 240,8)),
			7199 => std_logic_vector(to_unsigned( 115,8)),
			7200 => std_logic_vector(to_unsigned( 165,8)),
			7201 => std_logic_vector(to_unsigned( 187,8)),
			7202 => std_logic_vector(to_unsigned( 16,8)),
			7203 => std_logic_vector(to_unsigned( 172,8)),
			7204 => std_logic_vector(to_unsigned( 84,8)),
			7205 => std_logic_vector(to_unsigned( 104,8)),
			7206 => std_logic_vector(to_unsigned( 212,8)),
			7207 => std_logic_vector(to_unsigned( 19,8)),
			7208 => std_logic_vector(to_unsigned( 216,8)),
			7209 => std_logic_vector(to_unsigned( 34,8)),
			7210 => std_logic_vector(to_unsigned( 152,8)),
			7211 => std_logic_vector(to_unsigned( 11,8)),
			7212 => std_logic_vector(to_unsigned( 12,8)),
			7213 => std_logic_vector(to_unsigned( 154,8)),
			7214 => std_logic_vector(to_unsigned( 37,8)),
			7215 => std_logic_vector(to_unsigned( 207,8)),
			7216 => std_logic_vector(to_unsigned( 249,8)),
			7217 => std_logic_vector(to_unsigned( 177,8)),
			7218 => std_logic_vector(to_unsigned( 208,8)),
			7219 => std_logic_vector(to_unsigned( 72,8)),
			7220 => std_logic_vector(to_unsigned( 211,8)),
			7221 => std_logic_vector(to_unsigned( 132,8)),
			7222 => std_logic_vector(to_unsigned( 64,8)),
			7223 => std_logic_vector(to_unsigned( 16,8)),
			7224 => std_logic_vector(to_unsigned( 70,8)),
			7225 => std_logic_vector(to_unsigned( 158,8)),
			7226 => std_logic_vector(to_unsigned( 59,8)),
			7227 => std_logic_vector(to_unsigned( 110,8)),
			7228 => std_logic_vector(to_unsigned( 222,8)),
			7229 => std_logic_vector(to_unsigned( 218,8)),
			7230 => std_logic_vector(to_unsigned( 141,8)),
			7231 => std_logic_vector(to_unsigned( 65,8)),
			7232 => std_logic_vector(to_unsigned( 16,8)),
			7233 => std_logic_vector(to_unsigned( 186,8)),
			7234 => std_logic_vector(to_unsigned( 26,8)),
			7235 => std_logic_vector(to_unsigned( 146,8)),
			7236 => std_logic_vector(to_unsigned( 193,8)),
			7237 => std_logic_vector(to_unsigned( 253,8)),
			7238 => std_logic_vector(to_unsigned( 32,8)),
			7239 => std_logic_vector(to_unsigned( 225,8)),
			7240 => std_logic_vector(to_unsigned( 30,8)),
			7241 => std_logic_vector(to_unsigned( 58,8)),
			7242 => std_logic_vector(to_unsigned( 90,8)),
			7243 => std_logic_vector(to_unsigned( 56,8)),
			7244 => std_logic_vector(to_unsigned( 171,8)),
			7245 => std_logic_vector(to_unsigned( 159,8)),
			7246 => std_logic_vector(to_unsigned( 57,8)),
			7247 => std_logic_vector(to_unsigned( 164,8)),
			7248 => std_logic_vector(to_unsigned( 100,8)),
			7249 => std_logic_vector(to_unsigned( 115,8)),
			7250 => std_logic_vector(to_unsigned( 250,8)),
			7251 => std_logic_vector(to_unsigned( 12,8)),
			7252 => std_logic_vector(to_unsigned( 154,8)),
			7253 => std_logic_vector(to_unsigned( 238,8)),
			7254 => std_logic_vector(to_unsigned( 129,8)),
			7255 => std_logic_vector(to_unsigned( 248,8)),
			7256 => std_logic_vector(to_unsigned( 179,8)),
			7257 => std_logic_vector(to_unsigned( 131,8)),
			7258 => std_logic_vector(to_unsigned( 68,8)),
			7259 => std_logic_vector(to_unsigned( 77,8)),
			7260 => std_logic_vector(to_unsigned( 50,8)),
			7261 => std_logic_vector(to_unsigned( 83,8)),
			7262 => std_logic_vector(to_unsigned( 158,8)),
			7263 => std_logic_vector(to_unsigned( 164,8)),
			7264 => std_logic_vector(to_unsigned( 108,8)),
			7265 => std_logic_vector(to_unsigned( 44,8)),
			7266 => std_logic_vector(to_unsigned( 222,8)),
			7267 => std_logic_vector(to_unsigned( 221,8)),
			7268 => std_logic_vector(to_unsigned( 166,8)),
			7269 => std_logic_vector(to_unsigned( 242,8)),
			7270 => std_logic_vector(to_unsigned( 235,8)),
			7271 => std_logic_vector(to_unsigned( 56,8)),
			7272 => std_logic_vector(to_unsigned( 10,8)),
			7273 => std_logic_vector(to_unsigned( 29,8)),
			7274 => std_logic_vector(to_unsigned( 84,8)),
			7275 => std_logic_vector(to_unsigned( 205,8)),
			7276 => std_logic_vector(to_unsigned( 190,8)),
			7277 => std_logic_vector(to_unsigned( 224,8)),
			7278 => std_logic_vector(to_unsigned( 169,8)),
			7279 => std_logic_vector(to_unsigned( 97,8)),
			7280 => std_logic_vector(to_unsigned( 255,8)),
			7281 => std_logic_vector(to_unsigned( 141,8)),
			7282 => std_logic_vector(to_unsigned( 10,8)),
			7283 => std_logic_vector(to_unsigned( 182,8)),
			7284 => std_logic_vector(to_unsigned( 219,8)),
			7285 => std_logic_vector(to_unsigned( 6,8)),
			7286 => std_logic_vector(to_unsigned( 235,8)),
			7287 => std_logic_vector(to_unsigned( 162,8)),
			7288 => std_logic_vector(to_unsigned( 250,8)),
			7289 => std_logic_vector(to_unsigned( 9,8)),
			7290 => std_logic_vector(to_unsigned( 234,8)),
			7291 => std_logic_vector(to_unsigned( 40,8)),
			7292 => std_logic_vector(to_unsigned( 134,8)),
			7293 => std_logic_vector(to_unsigned( 92,8)),
			7294 => std_logic_vector(to_unsigned( 139,8)),
			7295 => std_logic_vector(to_unsigned( 52,8)),
			7296 => std_logic_vector(to_unsigned( 44,8)),
			7297 => std_logic_vector(to_unsigned( 223,8)),
			7298 => std_logic_vector(to_unsigned( 225,8)),
			7299 => std_logic_vector(to_unsigned( 188,8)),
			7300 => std_logic_vector(to_unsigned( 200,8)),
			7301 => std_logic_vector(to_unsigned( 112,8)),
			7302 => std_logic_vector(to_unsigned( 35,8)),
			7303 => std_logic_vector(to_unsigned( 140,8)),
			7304 => std_logic_vector(to_unsigned( 15,8)),
			7305 => std_logic_vector(to_unsigned( 5,8)),
			7306 => std_logic_vector(to_unsigned( 191,8)),
			7307 => std_logic_vector(to_unsigned( 104,8)),
			7308 => std_logic_vector(to_unsigned( 11,8)),
			7309 => std_logic_vector(to_unsigned( 128,8)),
			7310 => std_logic_vector(to_unsigned( 148,8)),
			7311 => std_logic_vector(to_unsigned( 8,8)),
			7312 => std_logic_vector(to_unsigned( 53,8)),
			7313 => std_logic_vector(to_unsigned( 220,8)),
			7314 => std_logic_vector(to_unsigned( 191,8)),
			7315 => std_logic_vector(to_unsigned( 67,8)),
			7316 => std_logic_vector(to_unsigned( 118,8)),
			7317 => std_logic_vector(to_unsigned( 94,8)),
			7318 => std_logic_vector(to_unsigned( 198,8)),
			7319 => std_logic_vector(to_unsigned( 18,8)),
			7320 => std_logic_vector(to_unsigned( 59,8)),
			7321 => std_logic_vector(to_unsigned( 241,8)),
			7322 => std_logic_vector(to_unsigned( 137,8)),
			7323 => std_logic_vector(to_unsigned( 130,8)),
			7324 => std_logic_vector(to_unsigned( 223,8)),
			7325 => std_logic_vector(to_unsigned( 90,8)),
			7326 => std_logic_vector(to_unsigned( 122,8)),
			7327 => std_logic_vector(to_unsigned( 252,8)),
			7328 => std_logic_vector(to_unsigned( 194,8)),
			7329 => std_logic_vector(to_unsigned( 132,8)),
			7330 => std_logic_vector(to_unsigned( 189,8)),
			7331 => std_logic_vector(to_unsigned( 204,8)),
			7332 => std_logic_vector(to_unsigned( 83,8)),
			7333 => std_logic_vector(to_unsigned( 228,8)),
			7334 => std_logic_vector(to_unsigned( 43,8)),
			7335 => std_logic_vector(to_unsigned( 147,8)),
			7336 => std_logic_vector(to_unsigned( 45,8)),
			7337 => std_logic_vector(to_unsigned( 8,8)),
			7338 => std_logic_vector(to_unsigned( 188,8)),
			7339 => std_logic_vector(to_unsigned( 111,8)),
			7340 => std_logic_vector(to_unsigned( 15,8)),
			7341 => std_logic_vector(to_unsigned( 72,8)),
			7342 => std_logic_vector(to_unsigned( 64,8)),
			7343 => std_logic_vector(to_unsigned( 172,8)),
			7344 => std_logic_vector(to_unsigned( 15,8)),
			7345 => std_logic_vector(to_unsigned( 95,8)),
			7346 => std_logic_vector(to_unsigned( 201,8)),
			7347 => std_logic_vector(to_unsigned( 120,8)),
			7348 => std_logic_vector(to_unsigned( 228,8)),
			7349 => std_logic_vector(to_unsigned( 194,8)),
			7350 => std_logic_vector(to_unsigned( 233,8)),
			7351 => std_logic_vector(to_unsigned( 76,8)),
			7352 => std_logic_vector(to_unsigned( 124,8)),
			7353 => std_logic_vector(to_unsigned( 150,8)),
			7354 => std_logic_vector(to_unsigned( 79,8)),
			7355 => std_logic_vector(to_unsigned( 159,8)),
			7356 => std_logic_vector(to_unsigned( 208,8)),
			7357 => std_logic_vector(to_unsigned( 211,8)),
			7358 => std_logic_vector(to_unsigned( 26,8)),
			7359 => std_logic_vector(to_unsigned( 29,8)),
			7360 => std_logic_vector(to_unsigned( 128,8)),
			7361 => std_logic_vector(to_unsigned( 37,8)),
			7362 => std_logic_vector(to_unsigned( 216,8)),
			7363 => std_logic_vector(to_unsigned( 246,8)),
			7364 => std_logic_vector(to_unsigned( 61,8)),
			7365 => std_logic_vector(to_unsigned( 102,8)),
			7366 => std_logic_vector(to_unsigned( 64,8)),
			7367 => std_logic_vector(to_unsigned( 71,8)),
			7368 => std_logic_vector(to_unsigned( 161,8)),
			7369 => std_logic_vector(to_unsigned( 248,8)),
			7370 => std_logic_vector(to_unsigned( 104,8)),
			7371 => std_logic_vector(to_unsigned( 232,8)),
			7372 => std_logic_vector(to_unsigned( 29,8)),
			7373 => std_logic_vector(to_unsigned( 72,8)),
			7374 => std_logic_vector(to_unsigned( 188,8)),
			7375 => std_logic_vector(to_unsigned( 8,8)),
			7376 => std_logic_vector(to_unsigned( 109,8)),
			7377 => std_logic_vector(to_unsigned( 155,8)),
			7378 => std_logic_vector(to_unsigned( 242,8)),
			7379 => std_logic_vector(to_unsigned( 179,8)),
			7380 => std_logic_vector(to_unsigned( 141,8)),
			7381 => std_logic_vector(to_unsigned( 170,8)),
			7382 => std_logic_vector(to_unsigned( 46,8)),
			7383 => std_logic_vector(to_unsigned( 31,8)),
			7384 => std_logic_vector(to_unsigned( 61,8)),
			7385 => std_logic_vector(to_unsigned( 21,8)),
			7386 => std_logic_vector(to_unsigned( 97,8)),
			7387 => std_logic_vector(to_unsigned( 80,8)),
			7388 => std_logic_vector(to_unsigned( 214,8)),
			7389 => std_logic_vector(to_unsigned( 241,8)),
			7390 => std_logic_vector(to_unsigned( 24,8)),
			7391 => std_logic_vector(to_unsigned( 150,8)),
			7392 => std_logic_vector(to_unsigned( 76,8)),
			7393 => std_logic_vector(to_unsigned( 7,8)),
			7394 => std_logic_vector(to_unsigned( 22,8)),
			7395 => std_logic_vector(to_unsigned( 144,8)),
			7396 => std_logic_vector(to_unsigned( 240,8)),
			7397 => std_logic_vector(to_unsigned( 220,8)),
			7398 => std_logic_vector(to_unsigned( 202,8)),
			7399 => std_logic_vector(to_unsigned( 238,8)),
			7400 => std_logic_vector(to_unsigned( 252,8)),
			7401 => std_logic_vector(to_unsigned( 74,8)),
			7402 => std_logic_vector(to_unsigned( 1,8)),
			7403 => std_logic_vector(to_unsigned( 54,8)),
			7404 => std_logic_vector(to_unsigned( 188,8)),
			7405 => std_logic_vector(to_unsigned( 212,8)),
			7406 => std_logic_vector(to_unsigned( 35,8)),
			7407 => std_logic_vector(to_unsigned( 191,8)),
			7408 => std_logic_vector(to_unsigned( 229,8)),
			7409 => std_logic_vector(to_unsigned( 201,8)),
			7410 => std_logic_vector(to_unsigned( 119,8)),
			7411 => std_logic_vector(to_unsigned( 203,8)),
			7412 => std_logic_vector(to_unsigned( 52,8)),
			7413 => std_logic_vector(to_unsigned( 229,8)),
			7414 => std_logic_vector(to_unsigned( 39,8)),
			7415 => std_logic_vector(to_unsigned( 112,8)),
			7416 => std_logic_vector(to_unsigned( 201,8)),
			7417 => std_logic_vector(to_unsigned( 101,8)),
			7418 => std_logic_vector(to_unsigned( 177,8)),
			7419 => std_logic_vector(to_unsigned( 191,8)),
			7420 => std_logic_vector(to_unsigned( 206,8)),
			7421 => std_logic_vector(to_unsigned( 28,8)),
			7422 => std_logic_vector(to_unsigned( 193,8)),
			7423 => std_logic_vector(to_unsigned( 208,8)),
			7424 => std_logic_vector(to_unsigned( 33,8)),
			7425 => std_logic_vector(to_unsigned( 147,8)),
			7426 => std_logic_vector(to_unsigned( 206,8)),
			7427 => std_logic_vector(to_unsigned( 98,8)),
			7428 => std_logic_vector(to_unsigned( 54,8)),
			7429 => std_logic_vector(to_unsigned( 54,8)),
			7430 => std_logic_vector(to_unsigned( 138,8)),
			7431 => std_logic_vector(to_unsigned( 225,8)),
			7432 => std_logic_vector(to_unsigned( 231,8)),
			7433 => std_logic_vector(to_unsigned( 21,8)),
			7434 => std_logic_vector(to_unsigned( 235,8)),
			7435 => std_logic_vector(to_unsigned( 134,8)),
			7436 => std_logic_vector(to_unsigned( 253,8)),
			7437 => std_logic_vector(to_unsigned( 126,8)),
			7438 => std_logic_vector(to_unsigned( 33,8)),
			7439 => std_logic_vector(to_unsigned( 170,8)),
			7440 => std_logic_vector(to_unsigned( 178,8)),
			7441 => std_logic_vector(to_unsigned( 187,8)),
			7442 => std_logic_vector(to_unsigned( 231,8)),
			7443 => std_logic_vector(to_unsigned( 173,8)),
			7444 => std_logic_vector(to_unsigned( 254,8)),
			7445 => std_logic_vector(to_unsigned( 37,8)),
			7446 => std_logic_vector(to_unsigned( 131,8)),
			7447 => std_logic_vector(to_unsigned( 107,8)),
			7448 => std_logic_vector(to_unsigned( 20,8)),
			7449 => std_logic_vector(to_unsigned( 253,8)),
			7450 => std_logic_vector(to_unsigned( 61,8)),
			7451 => std_logic_vector(to_unsigned( 175,8)),
			7452 => std_logic_vector(to_unsigned( 232,8)),
			7453 => std_logic_vector(to_unsigned( 152,8)),
			7454 => std_logic_vector(to_unsigned( 150,8)),
			7455 => std_logic_vector(to_unsigned( 208,8)),
			7456 => std_logic_vector(to_unsigned( 173,8)),
			7457 => std_logic_vector(to_unsigned( 204,8)),
			7458 => std_logic_vector(to_unsigned( 193,8)),
			7459 => std_logic_vector(to_unsigned( 31,8)),
			7460 => std_logic_vector(to_unsigned( 215,8)),
			7461 => std_logic_vector(to_unsigned( 239,8)),
			7462 => std_logic_vector(to_unsigned( 42,8)),
			7463 => std_logic_vector(to_unsigned( 68,8)),
			7464 => std_logic_vector(to_unsigned( 82,8)),
			7465 => std_logic_vector(to_unsigned( 221,8)),
			7466 => std_logic_vector(to_unsigned( 160,8)),
			7467 => std_logic_vector(to_unsigned( 227,8)),
			7468 => std_logic_vector(to_unsigned( 143,8)),
			7469 => std_logic_vector(to_unsigned( 34,8)),
			7470 => std_logic_vector(to_unsigned( 16,8)),
			7471 => std_logic_vector(to_unsigned( 54,8)),
			7472 => std_logic_vector(to_unsigned( 56,8)),
			7473 => std_logic_vector(to_unsigned( 11,8)),
			7474 => std_logic_vector(to_unsigned( 222,8)),
			7475 => std_logic_vector(to_unsigned( 113,8)),
			7476 => std_logic_vector(to_unsigned( 177,8)),
			7477 => std_logic_vector(to_unsigned( 99,8)),
			7478 => std_logic_vector(to_unsigned( 245,8)),
			7479 => std_logic_vector(to_unsigned( 103,8)),
			7480 => std_logic_vector(to_unsigned( 70,8)),
			7481 => std_logic_vector(to_unsigned( 72,8)),
			7482 => std_logic_vector(to_unsigned( 170,8)),
			7483 => std_logic_vector(to_unsigned( 113,8)),
			7484 => std_logic_vector(to_unsigned( 155,8)),
			7485 => std_logic_vector(to_unsigned( 178,8)),
			7486 => std_logic_vector(to_unsigned( 244,8)),
			7487 => std_logic_vector(to_unsigned( 28,8)),
			7488 => std_logic_vector(to_unsigned( 167,8)),
			7489 => std_logic_vector(to_unsigned( 90,8)),
			7490 => std_logic_vector(to_unsigned( 251,8)),
			7491 => std_logic_vector(to_unsigned( 62,8)),
			7492 => std_logic_vector(to_unsigned( 130,8)),
			7493 => std_logic_vector(to_unsigned( 132,8)),
			7494 => std_logic_vector(to_unsigned( 160,8)),
			7495 => std_logic_vector(to_unsigned( 173,8)),
			7496 => std_logic_vector(to_unsigned( 49,8)),
			7497 => std_logic_vector(to_unsigned( 69,8)),
			7498 => std_logic_vector(to_unsigned( 104,8)),
			7499 => std_logic_vector(to_unsigned( 0,8)),
			7500 => std_logic_vector(to_unsigned( 250,8)),
			7501 => std_logic_vector(to_unsigned( 65,8)),
			7502 => std_logic_vector(to_unsigned( 190,8)),
			7503 => std_logic_vector(to_unsigned( 40,8)),
			7504 => std_logic_vector(to_unsigned( 188,8)),
			7505 => std_logic_vector(to_unsigned( 112,8)),
			7506 => std_logic_vector(to_unsigned( 89,8)),
			7507 => std_logic_vector(to_unsigned( 68,8)),
			7508 => std_logic_vector(to_unsigned( 47,8)),
			7509 => std_logic_vector(to_unsigned( 21,8)),
			7510 => std_logic_vector(to_unsigned( 190,8)),
			7511 => std_logic_vector(to_unsigned( 170,8)),
			7512 => std_logic_vector(to_unsigned( 54,8)),
			7513 => std_logic_vector(to_unsigned( 35,8)),
			7514 => std_logic_vector(to_unsigned( 113,8)),
			7515 => std_logic_vector(to_unsigned( 135,8)),
			7516 => std_logic_vector(to_unsigned( 72,8)),
			7517 => std_logic_vector(to_unsigned( 189,8)),
			7518 => std_logic_vector(to_unsigned( 40,8)),
			7519 => std_logic_vector(to_unsigned( 23,8)),
			7520 => std_logic_vector(to_unsigned( 89,8)),
			7521 => std_logic_vector(to_unsigned( 254,8)),
			7522 => std_logic_vector(to_unsigned( 231,8)),
			7523 => std_logic_vector(to_unsigned( 142,8)),
			7524 => std_logic_vector(to_unsigned( 91,8)),
			7525 => std_logic_vector(to_unsigned( 109,8)),
			7526 => std_logic_vector(to_unsigned( 235,8)),
			7527 => std_logic_vector(to_unsigned( 111,8)),
			7528 => std_logic_vector(to_unsigned( 197,8)),
			7529 => std_logic_vector(to_unsigned( 65,8)),
			7530 => std_logic_vector(to_unsigned( 37,8)),
			7531 => std_logic_vector(to_unsigned( 129,8)),
			7532 => std_logic_vector(to_unsigned( 233,8)),
			7533 => std_logic_vector(to_unsigned( 24,8)),
			7534 => std_logic_vector(to_unsigned( 27,8)),
			7535 => std_logic_vector(to_unsigned( 79,8)),
			7536 => std_logic_vector(to_unsigned( 63,8)),
			7537 => std_logic_vector(to_unsigned( 21,8)),
			7538 => std_logic_vector(to_unsigned( 19,8)),
			7539 => std_logic_vector(to_unsigned( 29,8)),
			7540 => std_logic_vector(to_unsigned( 48,8)),
			7541 => std_logic_vector(to_unsigned( 212,8)),
			7542 => std_logic_vector(to_unsigned( 153,8)),
			7543 => std_logic_vector(to_unsigned( 57,8)),
			7544 => std_logic_vector(to_unsigned( 69,8)),
			7545 => std_logic_vector(to_unsigned( 247,8)),
			7546 => std_logic_vector(to_unsigned( 157,8)),
			7547 => std_logic_vector(to_unsigned( 98,8)),
			7548 => std_logic_vector(to_unsigned( 208,8)),
			7549 => std_logic_vector(to_unsigned( 109,8)),
			7550 => std_logic_vector(to_unsigned( 152,8)),
			7551 => std_logic_vector(to_unsigned( 149,8)),
			7552 => std_logic_vector(to_unsigned( 157,8)),
			7553 => std_logic_vector(to_unsigned( 135,8)),
			7554 => std_logic_vector(to_unsigned( 230,8)),
			7555 => std_logic_vector(to_unsigned( 185,8)),
			7556 => std_logic_vector(to_unsigned( 131,8)),
			7557 => std_logic_vector(to_unsigned( 71,8)),
			7558 => std_logic_vector(to_unsigned( 121,8)),
			7559 => std_logic_vector(to_unsigned( 184,8)),
			7560 => std_logic_vector(to_unsigned( 242,8)),
			7561 => std_logic_vector(to_unsigned( 149,8)),
			7562 => std_logic_vector(to_unsigned( 252,8)),
			7563 => std_logic_vector(to_unsigned( 101,8)),
			7564 => std_logic_vector(to_unsigned( 9,8)),
			7565 => std_logic_vector(to_unsigned( 72,8)),
			7566 => std_logic_vector(to_unsigned( 93,8)),
			7567 => std_logic_vector(to_unsigned( 2,8)),
			7568 => std_logic_vector(to_unsigned( 176,8)),
			7569 => std_logic_vector(to_unsigned( 140,8)),
			7570 => std_logic_vector(to_unsigned( 76,8)),
			7571 => std_logic_vector(to_unsigned( 236,8)),
			7572 => std_logic_vector(to_unsigned( 211,8)),
			7573 => std_logic_vector(to_unsigned( 111,8)),
			7574 => std_logic_vector(to_unsigned( 208,8)),
			7575 => std_logic_vector(to_unsigned( 62,8)),
			7576 => std_logic_vector(to_unsigned( 243,8)),
			7577 => std_logic_vector(to_unsigned( 42,8)),
			7578 => std_logic_vector(to_unsigned( 206,8)),
			7579 => std_logic_vector(to_unsigned( 174,8)),
			7580 => std_logic_vector(to_unsigned( 98,8)),
			7581 => std_logic_vector(to_unsigned( 198,8)),
			7582 => std_logic_vector(to_unsigned( 81,8)),
			7583 => std_logic_vector(to_unsigned( 176,8)),
			7584 => std_logic_vector(to_unsigned( 120,8)),
			7585 => std_logic_vector(to_unsigned( 171,8)),
			7586 => std_logic_vector(to_unsigned( 63,8)),
			7587 => std_logic_vector(to_unsigned( 64,8)),
			7588 => std_logic_vector(to_unsigned( 42,8)),
			7589 => std_logic_vector(to_unsigned( 202,8)),
			7590 => std_logic_vector(to_unsigned( 171,8)),
			7591 => std_logic_vector(to_unsigned( 159,8)),
			7592 => std_logic_vector(to_unsigned( 52,8)),
			7593 => std_logic_vector(to_unsigned( 181,8)),
			7594 => std_logic_vector(to_unsigned( 84,8)),
			7595 => std_logic_vector(to_unsigned( 184,8)),
			7596 => std_logic_vector(to_unsigned( 73,8)),
			7597 => std_logic_vector(to_unsigned( 175,8)),
			7598 => std_logic_vector(to_unsigned( 67,8)),
			7599 => std_logic_vector(to_unsigned( 52,8)),
			7600 => std_logic_vector(to_unsigned( 56,8)),
			7601 => std_logic_vector(to_unsigned( 49,8)),
			7602 => std_logic_vector(to_unsigned( 168,8)),
			7603 => std_logic_vector(to_unsigned( 35,8)),
			7604 => std_logic_vector(to_unsigned( 248,8)),
			7605 => std_logic_vector(to_unsigned( 224,8)),
			7606 => std_logic_vector(to_unsigned( 184,8)),
			7607 => std_logic_vector(to_unsigned( 152,8)),
			7608 => std_logic_vector(to_unsigned( 148,8)),
			7609 => std_logic_vector(to_unsigned( 1,8)),
			7610 => std_logic_vector(to_unsigned( 139,8)),
			7611 => std_logic_vector(to_unsigned( 56,8)),
			7612 => std_logic_vector(to_unsigned( 79,8)),
			7613 => std_logic_vector(to_unsigned( 139,8)),
			7614 => std_logic_vector(to_unsigned( 61,8)),
			7615 => std_logic_vector(to_unsigned( 73,8)),
			7616 => std_logic_vector(to_unsigned( 151,8)),
			7617 => std_logic_vector(to_unsigned( 218,8)),
			7618 => std_logic_vector(to_unsigned( 137,8)),
			7619 => std_logic_vector(to_unsigned( 42,8)),
			7620 => std_logic_vector(to_unsigned( 118,8)),
			7621 => std_logic_vector(to_unsigned( 115,8)),
			7622 => std_logic_vector(to_unsigned( 60,8)),
			7623 => std_logic_vector(to_unsigned( 110,8)),
			7624 => std_logic_vector(to_unsigned( 144,8)),
			7625 => std_logic_vector(to_unsigned( 174,8)),
			7626 => std_logic_vector(to_unsigned( 54,8)),
			7627 => std_logic_vector(to_unsigned( 158,8)),
			7628 => std_logic_vector(to_unsigned( 214,8)),
			7629 => std_logic_vector(to_unsigned( 87,8)),
			7630 => std_logic_vector(to_unsigned( 22,8)),
			7631 => std_logic_vector(to_unsigned( 116,8)),
			7632 => std_logic_vector(to_unsigned( 150,8)),
			7633 => std_logic_vector(to_unsigned( 237,8)),
			7634 => std_logic_vector(to_unsigned( 96,8)),
			7635 => std_logic_vector(to_unsigned( 19,8)),
			7636 => std_logic_vector(to_unsigned( 59,8)),
			7637 => std_logic_vector(to_unsigned( 121,8)),
			7638 => std_logic_vector(to_unsigned( 20,8)),
			7639 => std_logic_vector(to_unsigned( 122,8)),
			7640 => std_logic_vector(to_unsigned( 152,8)),
			7641 => std_logic_vector(to_unsigned( 99,8)),
			7642 => std_logic_vector(to_unsigned( 222,8)),
			7643 => std_logic_vector(to_unsigned( 68,8)),
			7644 => std_logic_vector(to_unsigned( 112,8)),
			7645 => std_logic_vector(to_unsigned( 171,8)),
			7646 => std_logic_vector(to_unsigned( 29,8)),
			7647 => std_logic_vector(to_unsigned( 207,8)),
			7648 => std_logic_vector(to_unsigned( 22,8)),
			7649 => std_logic_vector(to_unsigned( 77,8)),
			7650 => std_logic_vector(to_unsigned( 41,8)),
			7651 => std_logic_vector(to_unsigned( 189,8)),
			7652 => std_logic_vector(to_unsigned( 177,8)),
			7653 => std_logic_vector(to_unsigned( 240,8)),
			7654 => std_logic_vector(to_unsigned( 167,8)),
			7655 => std_logic_vector(to_unsigned( 22,8)),
			7656 => std_logic_vector(to_unsigned( 207,8)),
			7657 => std_logic_vector(to_unsigned( 94,8)),
			7658 => std_logic_vector(to_unsigned( 146,8)),
			7659 => std_logic_vector(to_unsigned( 25,8)),
			7660 => std_logic_vector(to_unsigned( 190,8)),
			7661 => std_logic_vector(to_unsigned( 24,8)),
			7662 => std_logic_vector(to_unsigned( 16,8)),
			7663 => std_logic_vector(to_unsigned( 49,8)),
			7664 => std_logic_vector(to_unsigned( 115,8)),
			7665 => std_logic_vector(to_unsigned( 180,8)),
			7666 => std_logic_vector(to_unsigned( 68,8)),
			7667 => std_logic_vector(to_unsigned( 214,8)),
			7668 => std_logic_vector(to_unsigned( 207,8)),
			7669 => std_logic_vector(to_unsigned( 248,8)),
			7670 => std_logic_vector(to_unsigned( 75,8)),
			7671 => std_logic_vector(to_unsigned( 52,8)),
			7672 => std_logic_vector(to_unsigned( 24,8)),
			7673 => std_logic_vector(to_unsigned( 227,8)),
			7674 => std_logic_vector(to_unsigned( 30,8)),
			7675 => std_logic_vector(to_unsigned( 171,8)),
			7676 => std_logic_vector(to_unsigned( 19,8)),
			7677 => std_logic_vector(to_unsigned( 167,8)),
			7678 => std_logic_vector(to_unsigned( 181,8)),
			7679 => std_logic_vector(to_unsigned( 224,8)),
			7680 => std_logic_vector(to_unsigned( 133,8)),
			7681 => std_logic_vector(to_unsigned( 248,8)),
			7682 => std_logic_vector(to_unsigned( 31,8)),
			7683 => std_logic_vector(to_unsigned( 201,8)),
			7684 => std_logic_vector(to_unsigned( 3,8)),
			7685 => std_logic_vector(to_unsigned( 90,8)),
			7686 => std_logic_vector(to_unsigned( 120,8)),
			7687 => std_logic_vector(to_unsigned( 231,8)),
			7688 => std_logic_vector(to_unsigned( 17,8)),
			7689 => std_logic_vector(to_unsigned( 64,8)),
			7690 => std_logic_vector(to_unsigned( 168,8)),
			7691 => std_logic_vector(to_unsigned( 180,8)),
			7692 => std_logic_vector(to_unsigned( 18,8)),
			7693 => std_logic_vector(to_unsigned( 82,8)),
			7694 => std_logic_vector(to_unsigned( 204,8)),
			7695 => std_logic_vector(to_unsigned( 68,8)),
			7696 => std_logic_vector(to_unsigned( 44,8)),
			7697 => std_logic_vector(to_unsigned( 124,8)),
			7698 => std_logic_vector(to_unsigned( 203,8)),
			7699 => std_logic_vector(to_unsigned( 233,8)),
			7700 => std_logic_vector(to_unsigned( 224,8)),
			7701 => std_logic_vector(to_unsigned( 239,8)),
			7702 => std_logic_vector(to_unsigned( 73,8)),
			7703 => std_logic_vector(to_unsigned( 156,8)),
			7704 => std_logic_vector(to_unsigned( 95,8)),
			7705 => std_logic_vector(to_unsigned( 157,8)),
			7706 => std_logic_vector(to_unsigned( 0,8)),
			7707 => std_logic_vector(to_unsigned( 129,8)),
			7708 => std_logic_vector(to_unsigned( 104,8)),
			7709 => std_logic_vector(to_unsigned( 11,8)),
			7710 => std_logic_vector(to_unsigned( 193,8)),
			7711 => std_logic_vector(to_unsigned( 199,8)),
			7712 => std_logic_vector(to_unsigned( 180,8)),
			7713 => std_logic_vector(to_unsigned( 116,8)),
			7714 => std_logic_vector(to_unsigned( 246,8)),
			7715 => std_logic_vector(to_unsigned( 2,8)),
			7716 => std_logic_vector(to_unsigned( 163,8)),
			7717 => std_logic_vector(to_unsigned( 96,8)),
			7718 => std_logic_vector(to_unsigned( 149,8)),
			7719 => std_logic_vector(to_unsigned( 64,8)),
			7720 => std_logic_vector(to_unsigned( 186,8)),
			7721 => std_logic_vector(to_unsigned( 166,8)),
			7722 => std_logic_vector(to_unsigned( 49,8)),
			7723 => std_logic_vector(to_unsigned( 116,8)),
			7724 => std_logic_vector(to_unsigned( 216,8)),
			7725 => std_logic_vector(to_unsigned( 104,8)),
			7726 => std_logic_vector(to_unsigned( 219,8)),
			7727 => std_logic_vector(to_unsigned( 88,8)),
			7728 => std_logic_vector(to_unsigned( 222,8)),
			7729 => std_logic_vector(to_unsigned( 165,8)),
			7730 => std_logic_vector(to_unsigned( 160,8)),
			7731 => std_logic_vector(to_unsigned( 254,8)),
			7732 => std_logic_vector(to_unsigned( 131,8)),
			7733 => std_logic_vector(to_unsigned( 40,8)),
			7734 => std_logic_vector(to_unsigned( 154,8)),
			7735 => std_logic_vector(to_unsigned( 139,8)),
			7736 => std_logic_vector(to_unsigned( 250,8)),
			7737 => std_logic_vector(to_unsigned( 117,8)),
			7738 => std_logic_vector(to_unsigned( 135,8)),
			7739 => std_logic_vector(to_unsigned( 3,8)),
			7740 => std_logic_vector(to_unsigned( 138,8)),
			7741 => std_logic_vector(to_unsigned( 237,8)),
			7742 => std_logic_vector(to_unsigned( 174,8)),
			7743 => std_logic_vector(to_unsigned( 179,8)),
			7744 => std_logic_vector(to_unsigned( 39,8)),
			7745 => std_logic_vector(to_unsigned( 121,8)),
			7746 => std_logic_vector(to_unsigned( 133,8)),
			7747 => std_logic_vector(to_unsigned( 64,8)),
			7748 => std_logic_vector(to_unsigned( 20,8)),
			7749 => std_logic_vector(to_unsigned( 74,8)),
			7750 => std_logic_vector(to_unsigned( 187,8)),
			7751 => std_logic_vector(to_unsigned( 87,8)),
			7752 => std_logic_vector(to_unsigned( 86,8)),
			7753 => std_logic_vector(to_unsigned( 200,8)),
			7754 => std_logic_vector(to_unsigned( 131,8)),
			7755 => std_logic_vector(to_unsigned( 64,8)),
			7756 => std_logic_vector(to_unsigned( 228,8)),
			7757 => std_logic_vector(to_unsigned( 185,8)),
			7758 => std_logic_vector(to_unsigned( 42,8)),
			7759 => std_logic_vector(to_unsigned( 54,8)),
			7760 => std_logic_vector(to_unsigned( 139,8)),
			7761 => std_logic_vector(to_unsigned( 218,8)),
			7762 => std_logic_vector(to_unsigned( 123,8)),
			7763 => std_logic_vector(to_unsigned( 91,8)),
			7764 => std_logic_vector(to_unsigned( 222,8)),
			7765 => std_logic_vector(to_unsigned( 52,8)),
			7766 => std_logic_vector(to_unsigned( 153,8)),
			7767 => std_logic_vector(to_unsigned( 40,8)),
			7768 => std_logic_vector(to_unsigned( 18,8)),
			7769 => std_logic_vector(to_unsigned( 209,8)),
			7770 => std_logic_vector(to_unsigned( 43,8)),
			7771 => std_logic_vector(to_unsigned( 33,8)),
			7772 => std_logic_vector(to_unsigned( 249,8)),
			7773 => std_logic_vector(to_unsigned( 22,8)),
			7774 => std_logic_vector(to_unsigned( 163,8)),
			7775 => std_logic_vector(to_unsigned( 12,8)),
			7776 => std_logic_vector(to_unsigned( 201,8)),
			7777 => std_logic_vector(to_unsigned( 64,8)),
			7778 => std_logic_vector(to_unsigned( 206,8)),
			7779 => std_logic_vector(to_unsigned( 249,8)),
			7780 => std_logic_vector(to_unsigned( 153,8)),
			7781 => std_logic_vector(to_unsigned( 126,8)),
			7782 => std_logic_vector(to_unsigned( 132,8)),
			7783 => std_logic_vector(to_unsigned( 255,8)),
			7784 => std_logic_vector(to_unsigned( 60,8)),
			7785 => std_logic_vector(to_unsigned( 156,8)),
			7786 => std_logic_vector(to_unsigned( 77,8)),
			7787 => std_logic_vector(to_unsigned( 190,8)),
			7788 => std_logic_vector(to_unsigned( 151,8)),
			7789 => std_logic_vector(to_unsigned( 111,8)),
			7790 => std_logic_vector(to_unsigned( 231,8)),
			7791 => std_logic_vector(to_unsigned( 251,8)),
			7792 => std_logic_vector(to_unsigned( 105,8)),
			7793 => std_logic_vector(to_unsigned( 176,8)),
			7794 => std_logic_vector(to_unsigned( 153,8)),
			7795 => std_logic_vector(to_unsigned( 146,8)),
			7796 => std_logic_vector(to_unsigned( 64,8)),
			7797 => std_logic_vector(to_unsigned( 195,8)),
			7798 => std_logic_vector(to_unsigned( 70,8)),
			7799 => std_logic_vector(to_unsigned( 229,8)),
			7800 => std_logic_vector(to_unsigned( 187,8)),
			7801 => std_logic_vector(to_unsigned( 62,8)),
			7802 => std_logic_vector(to_unsigned( 61,8)),
			7803 => std_logic_vector(to_unsigned( 44,8)),
			7804 => std_logic_vector(to_unsigned( 48,8)),
			7805 => std_logic_vector(to_unsigned( 127,8)),
			7806 => std_logic_vector(to_unsigned( 214,8)),
			7807 => std_logic_vector(to_unsigned( 167,8)),
			7808 => std_logic_vector(to_unsigned( 246,8)),
			7809 => std_logic_vector(to_unsigned( 0,8)),
			7810 => std_logic_vector(to_unsigned( 188,8)),
			7811 => std_logic_vector(to_unsigned( 118,8)),
			7812 => std_logic_vector(to_unsigned( 115,8)),
			7813 => std_logic_vector(to_unsigned( 220,8)),
			7814 => std_logic_vector(to_unsigned( 167,8)),
			7815 => std_logic_vector(to_unsigned( 90,8)),
			7816 => std_logic_vector(to_unsigned( 159,8)),
			7817 => std_logic_vector(to_unsigned( 199,8)),
			7818 => std_logic_vector(to_unsigned( 15,8)),
			7819 => std_logic_vector(to_unsigned( 90,8)),
			7820 => std_logic_vector(to_unsigned( 240,8)),
			7821 => std_logic_vector(to_unsigned( 147,8)),
			7822 => std_logic_vector(to_unsigned( 215,8)),
			7823 => std_logic_vector(to_unsigned( 2,8)),
			7824 => std_logic_vector(to_unsigned( 36,8)),
			7825 => std_logic_vector(to_unsigned( 106,8)),
			7826 => std_logic_vector(to_unsigned( 253,8)),
			7827 => std_logic_vector(to_unsigned( 18,8)),
			7828 => std_logic_vector(to_unsigned( 73,8)),
			7829 => std_logic_vector(to_unsigned( 44,8)),
			7830 => std_logic_vector(to_unsigned( 247,8)),
			7831 => std_logic_vector(to_unsigned( 197,8)),
			7832 => std_logic_vector(to_unsigned( 172,8)),
			7833 => std_logic_vector(to_unsigned( 220,8)),
			7834 => std_logic_vector(to_unsigned( 202,8)),
			7835 => std_logic_vector(to_unsigned( 123,8)),
			7836 => std_logic_vector(to_unsigned( 224,8)),
			7837 => std_logic_vector(to_unsigned( 241,8)),
			7838 => std_logic_vector(to_unsigned( 166,8)),
			7839 => std_logic_vector(to_unsigned( 36,8)),
			7840 => std_logic_vector(to_unsigned( 222,8)),
			7841 => std_logic_vector(to_unsigned( 139,8)),
			7842 => std_logic_vector(to_unsigned( 160,8)),
			7843 => std_logic_vector(to_unsigned( 0,8)),
			7844 => std_logic_vector(to_unsigned( 187,8)),
			7845 => std_logic_vector(to_unsigned( 190,8)),
			7846 => std_logic_vector(to_unsigned( 84,8)),
			7847 => std_logic_vector(to_unsigned( 124,8)),
			7848 => std_logic_vector(to_unsigned( 151,8)),
			7849 => std_logic_vector(to_unsigned( 90,8)),
			7850 => std_logic_vector(to_unsigned( 164,8)),
			7851 => std_logic_vector(to_unsigned( 103,8)),
			7852 => std_logic_vector(to_unsigned( 107,8)),
			7853 => std_logic_vector(to_unsigned( 222,8)),
			7854 => std_logic_vector(to_unsigned( 1,8)),
			7855 => std_logic_vector(to_unsigned( 245,8)),
			7856 => std_logic_vector(to_unsigned( 92,8)),
			7857 => std_logic_vector(to_unsigned( 60,8)),
			7858 => std_logic_vector(to_unsigned( 13,8)),
			7859 => std_logic_vector(to_unsigned( 216,8)),
			7860 => std_logic_vector(to_unsigned( 74,8)),
			7861 => std_logic_vector(to_unsigned( 53,8)),
			7862 => std_logic_vector(to_unsigned( 238,8)),
			7863 => std_logic_vector(to_unsigned( 23,8)),
			7864 => std_logic_vector(to_unsigned( 67,8)),
			7865 => std_logic_vector(to_unsigned( 157,8)),
			7866 => std_logic_vector(to_unsigned( 40,8)),
			7867 => std_logic_vector(to_unsigned( 108,8)),
			7868 => std_logic_vector(to_unsigned( 210,8)),
			7869 => std_logic_vector(to_unsigned( 63,8)),
			7870 => std_logic_vector(to_unsigned( 234,8)),
			7871 => std_logic_vector(to_unsigned( 76,8)),
			7872 => std_logic_vector(to_unsigned( 96,8)),
			7873 => std_logic_vector(to_unsigned( 134,8)),
			7874 => std_logic_vector(to_unsigned( 243,8)),
			7875 => std_logic_vector(to_unsigned( 213,8)),
			7876 => std_logic_vector(to_unsigned( 75,8)),
			7877 => std_logic_vector(to_unsigned( 217,8)),
			7878 => std_logic_vector(to_unsigned( 228,8)),
			7879 => std_logic_vector(to_unsigned( 42,8)),
			7880 => std_logic_vector(to_unsigned( 77,8)),
			7881 => std_logic_vector(to_unsigned( 163,8)),
			7882 => std_logic_vector(to_unsigned( 137,8)),
			7883 => std_logic_vector(to_unsigned( 108,8)),
			7884 => std_logic_vector(to_unsigned( 172,8)),
			7885 => std_logic_vector(to_unsigned( 59,8)),
			7886 => std_logic_vector(to_unsigned( 218,8)),
			7887 => std_logic_vector(to_unsigned( 170,8)),
			7888 => std_logic_vector(to_unsigned( 136,8)),
			7889 => std_logic_vector(to_unsigned( 176,8)),
			7890 => std_logic_vector(to_unsigned( 137,8)),
			7891 => std_logic_vector(to_unsigned( 120,8)),
			7892 => std_logic_vector(to_unsigned( 170,8)),
			7893 => std_logic_vector(to_unsigned( 75,8)),
			7894 => std_logic_vector(to_unsigned( 254,8)),
			7895 => std_logic_vector(to_unsigned( 221,8)),
			7896 => std_logic_vector(to_unsigned( 67,8)),
			7897 => std_logic_vector(to_unsigned( 171,8)),
			7898 => std_logic_vector(to_unsigned( 131,8)),
			7899 => std_logic_vector(to_unsigned( 176,8)),
			7900 => std_logic_vector(to_unsigned( 65,8)),
			7901 => std_logic_vector(to_unsigned( 145,8)),
			7902 => std_logic_vector(to_unsigned( 123,8)),
			7903 => std_logic_vector(to_unsigned( 208,8)),
			7904 => std_logic_vector(to_unsigned( 35,8)),
			7905 => std_logic_vector(to_unsigned( 213,8)),
			7906 => std_logic_vector(to_unsigned( 156,8)),
			7907 => std_logic_vector(to_unsigned( 199,8)),
			7908 => std_logic_vector(to_unsigned( 69,8)),
			7909 => std_logic_vector(to_unsigned( 36,8)),
			7910 => std_logic_vector(to_unsigned( 169,8)),
			7911 => std_logic_vector(to_unsigned( 218,8)),
			7912 => std_logic_vector(to_unsigned( 128,8)),
			7913 => std_logic_vector(to_unsigned( 156,8)),
			7914 => std_logic_vector(to_unsigned( 18,8)),
			7915 => std_logic_vector(to_unsigned( 126,8)),
			7916 => std_logic_vector(to_unsigned( 110,8)),
			7917 => std_logic_vector(to_unsigned( 207,8)),
			7918 => std_logic_vector(to_unsigned( 43,8)),
			7919 => std_logic_vector(to_unsigned( 11,8)),
			7920 => std_logic_vector(to_unsigned( 30,8)),
			7921 => std_logic_vector(to_unsigned( 206,8)),
			7922 => std_logic_vector(to_unsigned( 114,8)),
			7923 => std_logic_vector(to_unsigned( 222,8)),
			7924 => std_logic_vector(to_unsigned( 23,8)),
			7925 => std_logic_vector(to_unsigned( 169,8)),
			7926 => std_logic_vector(to_unsigned( 2,8)),
			7927 => std_logic_vector(to_unsigned( 218,8)),
			7928 => std_logic_vector(to_unsigned( 1,8)),
			7929 => std_logic_vector(to_unsigned( 89,8)),
			7930 => std_logic_vector(to_unsigned( 163,8)),
			7931 => std_logic_vector(to_unsigned( 162,8)),
			7932 => std_logic_vector(to_unsigned( 53,8)),
			7933 => std_logic_vector(to_unsigned( 131,8)),
			7934 => std_logic_vector(to_unsigned( 102,8)),
			7935 => std_logic_vector(to_unsigned( 182,8)),
			7936 => std_logic_vector(to_unsigned( 222,8)),
			7937 => std_logic_vector(to_unsigned( 28,8)),
			7938 => std_logic_vector(to_unsigned( 184,8)),
			7939 => std_logic_vector(to_unsigned( 189,8)),
			7940 => std_logic_vector(to_unsigned( 167,8)),
			7941 => std_logic_vector(to_unsigned( 186,8)),
			7942 => std_logic_vector(to_unsigned( 94,8)),
			7943 => std_logic_vector(to_unsigned( 53,8)),
			7944 => std_logic_vector(to_unsigned( 222,8)),
			7945 => std_logic_vector(to_unsigned( 32,8)),
			7946 => std_logic_vector(to_unsigned( 135,8)),
			7947 => std_logic_vector(to_unsigned( 126,8)),
			7948 => std_logic_vector(to_unsigned( 61,8)),
			7949 => std_logic_vector(to_unsigned( 238,8)),
			7950 => std_logic_vector(to_unsigned( 103,8)),
			7951 => std_logic_vector(to_unsigned( 68,8)),
			7952 => std_logic_vector(to_unsigned( 98,8)),
			7953 => std_logic_vector(to_unsigned( 76,8)),
			7954 => std_logic_vector(to_unsigned( 224,8)),
			7955 => std_logic_vector(to_unsigned( 167,8)),
			7956 => std_logic_vector(to_unsigned( 240,8)),
			7957 => std_logic_vector(to_unsigned( 0,8)),
			7958 => std_logic_vector(to_unsigned( 63,8)),
			7959 => std_logic_vector(to_unsigned( 34,8)),
			7960 => std_logic_vector(to_unsigned( 88,8)),
			7961 => std_logic_vector(to_unsigned( 226,8)),
			7962 => std_logic_vector(to_unsigned( 85,8)),
			7963 => std_logic_vector(to_unsigned( 134,8)),
			7964 => std_logic_vector(to_unsigned( 37,8)),
			7965 => std_logic_vector(to_unsigned( 157,8)),
			7966 => std_logic_vector(to_unsigned( 62,8)),
			7967 => std_logic_vector(to_unsigned( 34,8)),
			7968 => std_logic_vector(to_unsigned( 67,8)),
			7969 => std_logic_vector(to_unsigned( 117,8)),
			7970 => std_logic_vector(to_unsigned( 192,8)),
			7971 => std_logic_vector(to_unsigned( 132,8)),
			7972 => std_logic_vector(to_unsigned( 106,8)),
			7973 => std_logic_vector(to_unsigned( 88,8)),
			7974 => std_logic_vector(to_unsigned( 53,8)),
			7975 => std_logic_vector(to_unsigned( 193,8)),
			7976 => std_logic_vector(to_unsigned( 181,8)),
			7977 => std_logic_vector(to_unsigned( 165,8)),
			7978 => std_logic_vector(to_unsigned( 163,8)),
			7979 => std_logic_vector(to_unsigned( 46,8)),
			7980 => std_logic_vector(to_unsigned( 36,8)),
			7981 => std_logic_vector(to_unsigned( 227,8)),
			7982 => std_logic_vector(to_unsigned( 254,8)),
			7983 => std_logic_vector(to_unsigned( 240,8)),
			7984 => std_logic_vector(to_unsigned( 134,8)),
			7985 => std_logic_vector(to_unsigned( 27,8)),
			7986 => std_logic_vector(to_unsigned( 40,8)),
			7987 => std_logic_vector(to_unsigned( 113,8)),
			7988 => std_logic_vector(to_unsigned( 35,8)),
			7989 => std_logic_vector(to_unsigned( 173,8)),
			7990 => std_logic_vector(to_unsigned( 252,8)),
			7991 => std_logic_vector(to_unsigned( 241,8)),
			7992 => std_logic_vector(to_unsigned( 42,8)),
			7993 => std_logic_vector(to_unsigned( 212,8)),
			7994 => std_logic_vector(to_unsigned( 116,8)),
			7995 => std_logic_vector(to_unsigned( 98,8)),
			7996 => std_logic_vector(to_unsigned( 45,8)),
			7997 => std_logic_vector(to_unsigned( 64,8)),
			7998 => std_logic_vector(to_unsigned( 5,8)),
			7999 => std_logic_vector(to_unsigned( 84,8)),
			8000 => std_logic_vector(to_unsigned( 116,8)),
			8001 => std_logic_vector(to_unsigned( 39,8)),
			8002 => std_logic_vector(to_unsigned( 250,8)),
			8003 => std_logic_vector(to_unsigned( 4,8)),
			8004 => std_logic_vector(to_unsigned( 194,8)),
			8005 => std_logic_vector(to_unsigned( 115,8)),
			8006 => std_logic_vector(to_unsigned( 40,8)),
			8007 => std_logic_vector(to_unsigned( 89,8)),
			8008 => std_logic_vector(to_unsigned( 173,8)),
			8009 => std_logic_vector(to_unsigned( 28,8)),
			8010 => std_logic_vector(to_unsigned( 246,8)),
			8011 => std_logic_vector(to_unsigned( 99,8)),
			8012 => std_logic_vector(to_unsigned( 161,8)),
			8013 => std_logic_vector(to_unsigned( 29,8)),
			8014 => std_logic_vector(to_unsigned( 156,8)),
			8015 => std_logic_vector(to_unsigned( 89,8)),
			8016 => std_logic_vector(to_unsigned( 152,8)),
			8017 => std_logic_vector(to_unsigned( 201,8)),
			8018 => std_logic_vector(to_unsigned( 81,8)),
			8019 => std_logic_vector(to_unsigned( 27,8)),
			8020 => std_logic_vector(to_unsigned( 62,8)),
			8021 => std_logic_vector(to_unsigned( 148,8)),
			8022 => std_logic_vector(to_unsigned( 5,8)),
			8023 => std_logic_vector(to_unsigned( 193,8)),
			8024 => std_logic_vector(to_unsigned( 69,8)),
			8025 => std_logic_vector(to_unsigned( 246,8)),
			8026 => std_logic_vector(to_unsigned( 243,8)),
			8027 => std_logic_vector(to_unsigned( 85,8)),
			8028 => std_logic_vector(to_unsigned( 201,8)),
			8029 => std_logic_vector(to_unsigned( 132,8)),
			8030 => std_logic_vector(to_unsigned( 25,8)),
			8031 => std_logic_vector(to_unsigned( 97,8)),
			8032 => std_logic_vector(to_unsigned( 85,8)),
			8033 => std_logic_vector(to_unsigned( 207,8)),
			8034 => std_logic_vector(to_unsigned( 213,8)),
			8035 => std_logic_vector(to_unsigned( 237,8)),
			8036 => std_logic_vector(to_unsigned( 233,8)),
			8037 => std_logic_vector(to_unsigned( 150,8)),
			8038 => std_logic_vector(to_unsigned( 183,8)),
			8039 => std_logic_vector(to_unsigned( 165,8)),
			8040 => std_logic_vector(to_unsigned( 161,8)),
			8041 => std_logic_vector(to_unsigned( 179,8)),
			8042 => std_logic_vector(to_unsigned( 114,8)),
			8043 => std_logic_vector(to_unsigned( 22,8)),
			8044 => std_logic_vector(to_unsigned( 64,8)),
			8045 => std_logic_vector(to_unsigned( 163,8)),
			8046 => std_logic_vector(to_unsigned( 90,8)),
			8047 => std_logic_vector(to_unsigned( 172,8)),
			8048 => std_logic_vector(to_unsigned( 58,8)),
			8049 => std_logic_vector(to_unsigned( 41,8)),
			8050 => std_logic_vector(to_unsigned( 16,8)),
			8051 => std_logic_vector(to_unsigned( 162,8)),
			8052 => std_logic_vector(to_unsigned( 99,8)),
			8053 => std_logic_vector(to_unsigned( 101,8)),
			8054 => std_logic_vector(to_unsigned( 203,8)),
			8055 => std_logic_vector(to_unsigned( 142,8)),
			8056 => std_logic_vector(to_unsigned( 69,8)),
			8057 => std_logic_vector(to_unsigned( 67,8)),
			8058 => std_logic_vector(to_unsigned( 187,8)),
			8059 => std_logic_vector(to_unsigned( 145,8)),
			8060 => std_logic_vector(to_unsigned( 199,8)),
			8061 => std_logic_vector(to_unsigned( 145,8)),
			8062 => std_logic_vector(to_unsigned( 3,8)),
			8063 => std_logic_vector(to_unsigned( 30,8)),
			8064 => std_logic_vector(to_unsigned( 133,8)),
			8065 => std_logic_vector(to_unsigned( 6,8)),
			8066 => std_logic_vector(to_unsigned( 83,8)),
			8067 => std_logic_vector(to_unsigned( 150,8)),
			8068 => std_logic_vector(to_unsigned( 236,8)),
			8069 => std_logic_vector(to_unsigned( 206,8)),
			8070 => std_logic_vector(to_unsigned( 177,8)),
			8071 => std_logic_vector(to_unsigned( 112,8)),
			8072 => std_logic_vector(to_unsigned( 91,8)),
			8073 => std_logic_vector(to_unsigned( 190,8)),
			8074 => std_logic_vector(to_unsigned( 251,8)),
			8075 => std_logic_vector(to_unsigned( 198,8)),
			8076 => std_logic_vector(to_unsigned( 135,8)),
			8077 => std_logic_vector(to_unsigned( 36,8)),
			8078 => std_logic_vector(to_unsigned( 64,8)),
			8079 => std_logic_vector(to_unsigned( 119,8)),
			8080 => std_logic_vector(to_unsigned( 212,8)),
			8081 => std_logic_vector(to_unsigned( 83,8)),
			8082 => std_logic_vector(to_unsigned( 230,8)),
			8083 => std_logic_vector(to_unsigned( 253,8)),
			8084 => std_logic_vector(to_unsigned( 30,8)),
			8085 => std_logic_vector(to_unsigned( 33,8)),
			8086 => std_logic_vector(to_unsigned( 149,8)),
			8087 => std_logic_vector(to_unsigned( 179,8)),
			8088 => std_logic_vector(to_unsigned( 55,8)),
			8089 => std_logic_vector(to_unsigned( 210,8)),
			8090 => std_logic_vector(to_unsigned( 27,8)),
			8091 => std_logic_vector(to_unsigned( 19,8)),
			8092 => std_logic_vector(to_unsigned( 20,8)),
			8093 => std_logic_vector(to_unsigned( 146,8)),
			8094 => std_logic_vector(to_unsigned( 217,8)),
			8095 => std_logic_vector(to_unsigned( 239,8)),
			8096 => std_logic_vector(to_unsigned( 59,8)),
			8097 => std_logic_vector(to_unsigned( 106,8)),
			8098 => std_logic_vector(to_unsigned( 103,8)),
			8099 => std_logic_vector(to_unsigned( 220,8)),
			8100 => std_logic_vector(to_unsigned( 21,8)),
			8101 => std_logic_vector(to_unsigned( 132,8)),
			8102 => std_logic_vector(to_unsigned( 11,8)),
			8103 => std_logic_vector(to_unsigned( 185,8)),
			8104 => std_logic_vector(to_unsigned( 244,8)),
			8105 => std_logic_vector(to_unsigned( 94,8)),
			8106 => std_logic_vector(to_unsigned( 193,8)),
			8107 => std_logic_vector(to_unsigned( 21,8)),
			8108 => std_logic_vector(to_unsigned( 111,8)),
			8109 => std_logic_vector(to_unsigned( 255,8)),
			8110 => std_logic_vector(to_unsigned( 233,8)),
			8111 => std_logic_vector(to_unsigned( 23,8)),
			8112 => std_logic_vector(to_unsigned( 113,8)),
			8113 => std_logic_vector(to_unsigned( 51,8)),
			8114 => std_logic_vector(to_unsigned( 77,8)),
			8115 => std_logic_vector(to_unsigned( 248,8)),
			8116 => std_logic_vector(to_unsigned( 214,8)),
			8117 => std_logic_vector(to_unsigned( 3,8)),
			8118 => std_logic_vector(to_unsigned( 193,8)),
			8119 => std_logic_vector(to_unsigned( 71,8)),
			8120 => std_logic_vector(to_unsigned( 101,8)),
			8121 => std_logic_vector(to_unsigned( 208,8)),
			8122 => std_logic_vector(to_unsigned( 217,8)),
			8123 => std_logic_vector(to_unsigned( 20,8)),
			8124 => std_logic_vector(to_unsigned( 135,8)),
			8125 => std_logic_vector(to_unsigned( 174,8)),
			8126 => std_logic_vector(to_unsigned( 32,8)),
			8127 => std_logic_vector(to_unsigned( 189,8)),
			8128 => std_logic_vector(to_unsigned( 2,8)),
			8129 => std_logic_vector(to_unsigned( 200,8)),
			8130 => std_logic_vector(to_unsigned( 198,8)),
			8131 => std_logic_vector(to_unsigned( 5,8)),
			8132 => std_logic_vector(to_unsigned( 36,8)),
			8133 => std_logic_vector(to_unsigned( 24,8)),
			8134 => std_logic_vector(to_unsigned( 210,8)),
			8135 => std_logic_vector(to_unsigned( 103,8)),
			8136 => std_logic_vector(to_unsigned( 8,8)),
			8137 => std_logic_vector(to_unsigned( 141,8)),
			8138 => std_logic_vector(to_unsigned( 119,8)),
			8139 => std_logic_vector(to_unsigned( 186,8)),
			8140 => std_logic_vector(to_unsigned( 35,8)),
			8141 => std_logic_vector(to_unsigned( 148,8)),
			8142 => std_logic_vector(to_unsigned( 37,8)),
			8143 => std_logic_vector(to_unsigned( 68,8)),
			8144 => std_logic_vector(to_unsigned( 254,8)),
			8145 => std_logic_vector(to_unsigned( 251,8)),
			8146 => std_logic_vector(to_unsigned( 19,8)),
			8147 => std_logic_vector(to_unsigned( 96,8)),
			8148 => std_logic_vector(to_unsigned( 230,8)),
			8149 => std_logic_vector(to_unsigned( 166,8)),
			8150 => std_logic_vector(to_unsigned( 193,8)),
			8151 => std_logic_vector(to_unsigned( 162,8)),
			8152 => std_logic_vector(to_unsigned( 93,8)),
			8153 => std_logic_vector(to_unsigned( 7,8)),
			8154 => std_logic_vector(to_unsigned( 95,8)),
			8155 => std_logic_vector(to_unsigned( 174,8)),
			8156 => std_logic_vector(to_unsigned( 1,8)),
			8157 => std_logic_vector(to_unsigned( 208,8)),
			8158 => std_logic_vector(to_unsigned( 181,8)),
			8159 => std_logic_vector(to_unsigned( 216,8)),
			8160 => std_logic_vector(to_unsigned( 200,8)),
			8161 => std_logic_vector(to_unsigned( 137,8)),
			8162 => std_logic_vector(to_unsigned( 89,8)),
			8163 => std_logic_vector(to_unsigned( 74,8)),
			8164 => std_logic_vector(to_unsigned( 148,8)),
			8165 => std_logic_vector(to_unsigned( 163,8)),
			8166 => std_logic_vector(to_unsigned( 148,8)),
			8167 => std_logic_vector(to_unsigned( 39,8)),
			8168 => std_logic_vector(to_unsigned( 14,8)),
			8169 => std_logic_vector(to_unsigned( 86,8)),
			8170 => std_logic_vector(to_unsigned( 204,8)),
			8171 => std_logic_vector(to_unsigned( 105,8)),
			8172 => std_logic_vector(to_unsigned( 34,8)),
			8173 => std_logic_vector(to_unsigned( 18,8)),
			8174 => std_logic_vector(to_unsigned( 167,8)),
			8175 => std_logic_vector(to_unsigned( 15,8)),
			8176 => std_logic_vector(to_unsigned( 111,8)),
			8177 => std_logic_vector(to_unsigned( 20,8)),
			8178 => std_logic_vector(to_unsigned( 235,8)),
			8179 => std_logic_vector(to_unsigned( 8,8)),
			8180 => std_logic_vector(to_unsigned( 113,8)),
			8181 => std_logic_vector(to_unsigned( 204,8)),
			8182 => std_logic_vector(to_unsigned( 29,8)),
			8183 => std_logic_vector(to_unsigned( 156,8)),
			8184 => std_logic_vector(to_unsigned( 120,8)),
			8185 => std_logic_vector(to_unsigned( 19,8)),
			8186 => std_logic_vector(to_unsigned( 16,8)),
			8187 => std_logic_vector(to_unsigned( 196,8)),
			8188 => std_logic_vector(to_unsigned( 169,8)),
			8189 => std_logic_vector(to_unsigned( 194,8)),
			8190 => std_logic_vector(to_unsigned( 82,8)),
			8191 => std_logic_vector(to_unsigned( 29,8)),
			8192 => std_logic_vector(to_unsigned( 181,8)),
			8193 => std_logic_vector(to_unsigned( 121,8)),
			8194 => std_logic_vector(to_unsigned( 9,8)),
			8195 => std_logic_vector(to_unsigned( 112,8)),
			8196 => std_logic_vector(to_unsigned( 176,8)),
			8197 => std_logic_vector(to_unsigned( 6,8)),
			8198 => std_logic_vector(to_unsigned( 203,8)),
			8199 => std_logic_vector(to_unsigned( 16,8)),
			8200 => std_logic_vector(to_unsigned( 238,8)),
			8201 => std_logic_vector(to_unsigned( 39,8)),
			8202 => std_logic_vector(to_unsigned( 21,8)),
			8203 => std_logic_vector(to_unsigned( 165,8)),
			8204 => std_logic_vector(to_unsigned( 240,8)),
			8205 => std_logic_vector(to_unsigned( 34,8)),
			8206 => std_logic_vector(to_unsigned( 235,8)),
			8207 => std_logic_vector(to_unsigned( 164,8)),
			8208 => std_logic_vector(to_unsigned( 205,8)),
			8209 => std_logic_vector(to_unsigned( 215,8)),
			8210 => std_logic_vector(to_unsigned( 87,8)),
			8211 => std_logic_vector(to_unsigned( 90,8)),
			8212 => std_logic_vector(to_unsigned( 147,8)),
			8213 => std_logic_vector(to_unsigned( 233,8)),
			8214 => std_logic_vector(to_unsigned( 128,8)),
			8215 => std_logic_vector(to_unsigned( 189,8)),
			8216 => std_logic_vector(to_unsigned( 106,8)),
			8217 => std_logic_vector(to_unsigned( 160,8)),
			8218 => std_logic_vector(to_unsigned( 221,8)),
			8219 => std_logic_vector(to_unsigned( 43,8)),
			8220 => std_logic_vector(to_unsigned( 23,8)),
			8221 => std_logic_vector(to_unsigned( 193,8)),
			8222 => std_logic_vector(to_unsigned( 7,8)),
			8223 => std_logic_vector(to_unsigned( 96,8)),
			8224 => std_logic_vector(to_unsigned( 236,8)),
			8225 => std_logic_vector(to_unsigned( 148,8)),
			8226 => std_logic_vector(to_unsigned( 152,8)),
			8227 => std_logic_vector(to_unsigned( 148,8)),
			8228 => std_logic_vector(to_unsigned( 211,8)),
			8229 => std_logic_vector(to_unsigned( 7,8)),
			8230 => std_logic_vector(to_unsigned( 208,8)),
			8231 => std_logic_vector(to_unsigned( 52,8)),
			8232 => std_logic_vector(to_unsigned( 11,8)),
			8233 => std_logic_vector(to_unsigned( 181,8)),
			8234 => std_logic_vector(to_unsigned( 189,8)),
			8235 => std_logic_vector(to_unsigned( 165,8)),
			8236 => std_logic_vector(to_unsigned( 214,8)),
			8237 => std_logic_vector(to_unsigned( 214,8)),
			8238 => std_logic_vector(to_unsigned( 192,8)),
			8239 => std_logic_vector(to_unsigned( 176,8)),
			8240 => std_logic_vector(to_unsigned( 61,8)),
			8241 => std_logic_vector(to_unsigned( 140,8)),
			8242 => std_logic_vector(to_unsigned( 56,8)),
			8243 => std_logic_vector(to_unsigned( 0,8)),
			8244 => std_logic_vector(to_unsigned( 132,8)),
			8245 => std_logic_vector(to_unsigned( 23,8)),
			8246 => std_logic_vector(to_unsigned( 217,8)),
			8247 => std_logic_vector(to_unsigned( 241,8)),
			8248 => std_logic_vector(to_unsigned( 203,8)),
			8249 => std_logic_vector(to_unsigned( 78,8)),
			8250 => std_logic_vector(to_unsigned( 15,8)),
			8251 => std_logic_vector(to_unsigned( 36,8)),
			8252 => std_logic_vector(to_unsigned( 118,8)),
			8253 => std_logic_vector(to_unsigned( 255,8)),
			8254 => std_logic_vector(to_unsigned( 76,8)),
			8255 => std_logic_vector(to_unsigned( 188,8)),
			8256 => std_logic_vector(to_unsigned( 134,8)),
			8257 => std_logic_vector(to_unsigned( 145,8)),
			8258 => std_logic_vector(to_unsigned( 15,8)),
			8259 => std_logic_vector(to_unsigned( 22,8)),
			8260 => std_logic_vector(to_unsigned( 213,8)),
			8261 => std_logic_vector(to_unsigned( 92,8)),
			8262 => std_logic_vector(to_unsigned( 123,8)),
			8263 => std_logic_vector(to_unsigned( 203,8)),
			8264 => std_logic_vector(to_unsigned( 101,8)),
			8265 => std_logic_vector(to_unsigned( 76,8)),
			8266 => std_logic_vector(to_unsigned( 166,8)),
			8267 => std_logic_vector(to_unsigned( 81,8)),
			8268 => std_logic_vector(to_unsigned( 140,8)),
			8269 => std_logic_vector(to_unsigned( 208,8)),
			8270 => std_logic_vector(to_unsigned( 175,8)),
			8271 => std_logic_vector(to_unsigned( 72,8)),
			8272 => std_logic_vector(to_unsigned( 75,8)),
			8273 => std_logic_vector(to_unsigned( 192,8)),
			8274 => std_logic_vector(to_unsigned( 64,8)),
			8275 => std_logic_vector(to_unsigned( 238,8)),
			8276 => std_logic_vector(to_unsigned( 109,8)),
			8277 => std_logic_vector(to_unsigned( 174,8)),
			8278 => std_logic_vector(to_unsigned( 129,8)),
			8279 => std_logic_vector(to_unsigned( 73,8)),
			8280 => std_logic_vector(to_unsigned( 62,8)),
			8281 => std_logic_vector(to_unsigned( 241,8)),
			8282 => std_logic_vector(to_unsigned( 49,8)),
			8283 => std_logic_vector(to_unsigned( 2,8)),
			8284 => std_logic_vector(to_unsigned( 19,8)),
			8285 => std_logic_vector(to_unsigned( 106,8)),
			8286 => std_logic_vector(to_unsigned( 255,8)),
			8287 => std_logic_vector(to_unsigned( 143,8)),
			8288 => std_logic_vector(to_unsigned( 56,8)),
			8289 => std_logic_vector(to_unsigned( 45,8)),
			8290 => std_logic_vector(to_unsigned( 175,8)),
			8291 => std_logic_vector(to_unsigned( 242,8)),
			8292 => std_logic_vector(to_unsigned( 169,8)),
			8293 => std_logic_vector(to_unsigned( 6,8)),
			8294 => std_logic_vector(to_unsigned( 125,8)),
			8295 => std_logic_vector(to_unsigned( 57,8)),
			8296 => std_logic_vector(to_unsigned( 109,8)),
			8297 => std_logic_vector(to_unsigned( 2,8)),
			8298 => std_logic_vector(to_unsigned( 100,8)),
			8299 => std_logic_vector(to_unsigned( 228,8)),
			8300 => std_logic_vector(to_unsigned( 234,8)),
			8301 => std_logic_vector(to_unsigned( 95,8)),
			8302 => std_logic_vector(to_unsigned( 212,8)),
			8303 => std_logic_vector(to_unsigned( 85,8)),
			8304 => std_logic_vector(to_unsigned( 55,8)),
			8305 => std_logic_vector(to_unsigned( 175,8)),
			8306 => std_logic_vector(to_unsigned( 95,8)),
			8307 => std_logic_vector(to_unsigned( 185,8)),
			8308 => std_logic_vector(to_unsigned( 191,8)),
			8309 => std_logic_vector(to_unsigned( 114,8)),
			8310 => std_logic_vector(to_unsigned( 90,8)),
			8311 => std_logic_vector(to_unsigned( 8,8)),
			8312 => std_logic_vector(to_unsigned( 92,8)),
			8313 => std_logic_vector(to_unsigned( 245,8)),
			8314 => std_logic_vector(to_unsigned( 185,8)),
			8315 => std_logic_vector(to_unsigned( 224,8)),
			8316 => std_logic_vector(to_unsigned( 91,8)),
			8317 => std_logic_vector(to_unsigned( 55,8)),
			8318 => std_logic_vector(to_unsigned( 226,8)),
			8319 => std_logic_vector(to_unsigned( 73,8)),
			8320 => std_logic_vector(to_unsigned( 132,8)),
			8321 => std_logic_vector(to_unsigned( 147,8)),
			8322 => std_logic_vector(to_unsigned( 119,8)),
			8323 => std_logic_vector(to_unsigned( 203,8)),
			8324 => std_logic_vector(to_unsigned( 76,8)),
			8325 => std_logic_vector(to_unsigned( 24,8)),
			8326 => std_logic_vector(to_unsigned( 118,8)),
			8327 => std_logic_vector(to_unsigned( 71,8)),
			8328 => std_logic_vector(to_unsigned( 114,8)),
			8329 => std_logic_vector(to_unsigned( 202,8)),
			8330 => std_logic_vector(to_unsigned( 27,8)),
			8331 => std_logic_vector(to_unsigned( 221,8)),
			8332 => std_logic_vector(to_unsigned( 170,8)),
			8333 => std_logic_vector(to_unsigned( 102,8)),
			8334 => std_logic_vector(to_unsigned( 117,8)),
			8335 => std_logic_vector(to_unsigned( 90,8)),
			8336 => std_logic_vector(to_unsigned( 83,8)),
			8337 => std_logic_vector(to_unsigned( 151,8)),
			8338 => std_logic_vector(to_unsigned( 236,8)),
			8339 => std_logic_vector(to_unsigned( 92,8)),
			8340 => std_logic_vector(to_unsigned( 201,8)),
			8341 => std_logic_vector(to_unsigned( 66,8)),
			8342 => std_logic_vector(to_unsigned( 218,8)),
			8343 => std_logic_vector(to_unsigned( 75,8)),
			8344 => std_logic_vector(to_unsigned( 154,8)),
			8345 => std_logic_vector(to_unsigned( 110,8)),
			8346 => std_logic_vector(to_unsigned( 50,8)),
			8347 => std_logic_vector(to_unsigned( 148,8)),
			8348 => std_logic_vector(to_unsigned( 32,8)),
			8349 => std_logic_vector(to_unsigned( 151,8)),
			8350 => std_logic_vector(to_unsigned( 198,8)),
			8351 => std_logic_vector(to_unsigned( 76,8)),
			8352 => std_logic_vector(to_unsigned( 125,8)),
			8353 => std_logic_vector(to_unsigned( 236,8)),
			8354 => std_logic_vector(to_unsigned( 249,8)),
			8355 => std_logic_vector(to_unsigned( 124,8)),
			8356 => std_logic_vector(to_unsigned( 122,8)),
			8357 => std_logic_vector(to_unsigned( 73,8)),
			8358 => std_logic_vector(to_unsigned( 171,8)),
			8359 => std_logic_vector(to_unsigned( 144,8)),
			8360 => std_logic_vector(to_unsigned( 245,8)),
			8361 => std_logic_vector(to_unsigned( 3,8)),
			8362 => std_logic_vector(to_unsigned( 25,8)),
			8363 => std_logic_vector(to_unsigned( 70,8)),
			8364 => std_logic_vector(to_unsigned( 206,8)),
			8365 => std_logic_vector(to_unsigned( 185,8)),
			8366 => std_logic_vector(to_unsigned( 201,8)),
			8367 => std_logic_vector(to_unsigned( 254,8)),
			8368 => std_logic_vector(to_unsigned( 29,8)),
			8369 => std_logic_vector(to_unsigned( 213,8)),
			8370 => std_logic_vector(to_unsigned( 201,8)),
			8371 => std_logic_vector(to_unsigned( 231,8)),
			8372 => std_logic_vector(to_unsigned( 95,8)),
			8373 => std_logic_vector(to_unsigned( 43,8)),
			8374 => std_logic_vector(to_unsigned( 225,8)),
			8375 => std_logic_vector(to_unsigned( 243,8)),
			8376 => std_logic_vector(to_unsigned( 193,8)),
			8377 => std_logic_vector(to_unsigned( 23,8)),
			8378 => std_logic_vector(to_unsigned( 196,8)),
			8379 => std_logic_vector(to_unsigned( 234,8)),
			8380 => std_logic_vector(to_unsigned( 123,8)),
			8381 => std_logic_vector(to_unsigned( 206,8)),
			8382 => std_logic_vector(to_unsigned( 240,8)),
			8383 => std_logic_vector(to_unsigned( 220,8)),
			8384 => std_logic_vector(to_unsigned( 246,8)),
			8385 => std_logic_vector(to_unsigned( 115,8)),
			8386 => std_logic_vector(to_unsigned( 233,8)),
			8387 => std_logic_vector(to_unsigned( 163,8)),
			8388 => std_logic_vector(to_unsigned( 59,8)),
			8389 => std_logic_vector(to_unsigned( 145,8)),
			8390 => std_logic_vector(to_unsigned( 9,8)),
			8391 => std_logic_vector(to_unsigned( 49,8)),
			8392 => std_logic_vector(to_unsigned( 77,8)),
			8393 => std_logic_vector(to_unsigned( 237,8)),
			8394 => std_logic_vector(to_unsigned( 199,8)),
			8395 => std_logic_vector(to_unsigned( 17,8)),
			8396 => std_logic_vector(to_unsigned( 181,8)),
			8397 => std_logic_vector(to_unsigned( 162,8)),
			8398 => std_logic_vector(to_unsigned( 40,8)),
			8399 => std_logic_vector(to_unsigned( 29,8)),
			8400 => std_logic_vector(to_unsigned( 245,8)),
			8401 => std_logic_vector(to_unsigned( 20,8)),
			8402 => std_logic_vector(to_unsigned( 213,8)),
			8403 => std_logic_vector(to_unsigned( 132,8)),
			8404 => std_logic_vector(to_unsigned( 52,8)),
			8405 => std_logic_vector(to_unsigned( 219,8)),
			8406 => std_logic_vector(to_unsigned( 90,8)),
			8407 => std_logic_vector(to_unsigned( 22,8)),
			8408 => std_logic_vector(to_unsigned( 161,8)),
			8409 => std_logic_vector(to_unsigned( 53,8)),
			8410 => std_logic_vector(to_unsigned( 33,8)),
			8411 => std_logic_vector(to_unsigned( 196,8)),
			8412 => std_logic_vector(to_unsigned( 104,8)),
			8413 => std_logic_vector(to_unsigned( 108,8)),
			8414 => std_logic_vector(to_unsigned( 201,8)),
			8415 => std_logic_vector(to_unsigned( 103,8)),
			8416 => std_logic_vector(to_unsigned( 49,8)),
			8417 => std_logic_vector(to_unsigned( 71,8)),
			8418 => std_logic_vector(to_unsigned( 223,8)),
			8419 => std_logic_vector(to_unsigned( 69,8)),
			8420 => std_logic_vector(to_unsigned( 110,8)),
			8421 => std_logic_vector(to_unsigned( 61,8)),
			8422 => std_logic_vector(to_unsigned( 76,8)),
			8423 => std_logic_vector(to_unsigned( 21,8)),
			8424 => std_logic_vector(to_unsigned( 41,8)),
			8425 => std_logic_vector(to_unsigned( 241,8)),
			8426 => std_logic_vector(to_unsigned( 240,8)),
			8427 => std_logic_vector(to_unsigned( 186,8)),
			8428 => std_logic_vector(to_unsigned( 160,8)),
			8429 => std_logic_vector(to_unsigned( 152,8)),
			8430 => std_logic_vector(to_unsigned( 170,8)),
			8431 => std_logic_vector(to_unsigned( 249,8)),
			8432 => std_logic_vector(to_unsigned( 161,8)),
			8433 => std_logic_vector(to_unsigned( 117,8)),
			8434 => std_logic_vector(to_unsigned( 220,8)),
			8435 => std_logic_vector(to_unsigned( 54,8)),
			8436 => std_logic_vector(to_unsigned( 94,8)),
			8437 => std_logic_vector(to_unsigned( 149,8)),
			8438 => std_logic_vector(to_unsigned( 28,8)),
			8439 => std_logic_vector(to_unsigned( 103,8)),
			8440 => std_logic_vector(to_unsigned( 86,8)),
			8441 => std_logic_vector(to_unsigned( 200,8)),
			8442 => std_logic_vector(to_unsigned( 224,8)),
			8443 => std_logic_vector(to_unsigned( 202,8)),
			8444 => std_logic_vector(to_unsigned( 133,8)),
			8445 => std_logic_vector(to_unsigned( 188,8)),
			8446 => std_logic_vector(to_unsigned( 237,8)),
			8447 => std_logic_vector(to_unsigned( 236,8)),
			8448 => std_logic_vector(to_unsigned( 134,8)),
			8449 => std_logic_vector(to_unsigned( 120,8)),
			8450 => std_logic_vector(to_unsigned( 34,8)),
			8451 => std_logic_vector(to_unsigned( 203,8)),
			8452 => std_logic_vector(to_unsigned( 161,8)),
			8453 => std_logic_vector(to_unsigned( 36,8)),
			8454 => std_logic_vector(to_unsigned( 23,8)),
			8455 => std_logic_vector(to_unsigned( 120,8)),
			8456 => std_logic_vector(to_unsigned( 92,8)),
			8457 => std_logic_vector(to_unsigned( 174,8)),
			8458 => std_logic_vector(to_unsigned( 27,8)),
			8459 => std_logic_vector(to_unsigned( 177,8)),
			8460 => std_logic_vector(to_unsigned( 144,8)),
			8461 => std_logic_vector(to_unsigned( 153,8)),
			8462 => std_logic_vector(to_unsigned( 249,8)),
			8463 => std_logic_vector(to_unsigned( 247,8)),
			8464 => std_logic_vector(to_unsigned( 188,8)),
			8465 => std_logic_vector(to_unsigned( 195,8)),
			8466 => std_logic_vector(to_unsigned( 42,8)),
			8467 => std_logic_vector(to_unsigned( 237,8)),
			8468 => std_logic_vector(to_unsigned( 173,8)),
			8469 => std_logic_vector(to_unsigned( 142,8)),
			8470 => std_logic_vector(to_unsigned( 78,8)),
			8471 => std_logic_vector(to_unsigned( 152,8)),
			8472 => std_logic_vector(to_unsigned( 45,8)),
			8473 => std_logic_vector(to_unsigned( 159,8)),
			8474 => std_logic_vector(to_unsigned( 161,8)),
			8475 => std_logic_vector(to_unsigned( 103,8)),
			8476 => std_logic_vector(to_unsigned( 9,8)),
			8477 => std_logic_vector(to_unsigned( 249,8)),
			8478 => std_logic_vector(to_unsigned( 84,8)),
			8479 => std_logic_vector(to_unsigned( 57,8)),
			8480 => std_logic_vector(to_unsigned( 20,8)),
			8481 => std_logic_vector(to_unsigned( 54,8)),
			8482 => std_logic_vector(to_unsigned( 44,8)),
			8483 => std_logic_vector(to_unsigned( 52,8)),
			8484 => std_logic_vector(to_unsigned( 3,8)),
			8485 => std_logic_vector(to_unsigned( 154,8)),
			8486 => std_logic_vector(to_unsigned( 102,8)),
			8487 => std_logic_vector(to_unsigned( 141,8)),
			8488 => std_logic_vector(to_unsigned( 167,8)),
			8489 => std_logic_vector(to_unsigned( 158,8)),
			8490 => std_logic_vector(to_unsigned( 75,8)),
			8491 => std_logic_vector(to_unsigned( 74,8)),
			8492 => std_logic_vector(to_unsigned( 121,8)),
			8493 => std_logic_vector(to_unsigned( 144,8)),
			8494 => std_logic_vector(to_unsigned( 12,8)),
			8495 => std_logic_vector(to_unsigned( 182,8)),
			8496 => std_logic_vector(to_unsigned( 197,8)),
			8497 => std_logic_vector(to_unsigned( 82,8)),
			8498 => std_logic_vector(to_unsigned( 102,8)),
			8499 => std_logic_vector(to_unsigned( 143,8)),
			8500 => std_logic_vector(to_unsigned( 184,8)),
			8501 => std_logic_vector(to_unsigned( 15,8)),
			8502 => std_logic_vector(to_unsigned( 69,8)),
			8503 => std_logic_vector(to_unsigned( 133,8)),
			8504 => std_logic_vector(to_unsigned( 251,8)),
			8505 => std_logic_vector(to_unsigned( 116,8)),
			8506 => std_logic_vector(to_unsigned( 187,8)),
			8507 => std_logic_vector(to_unsigned( 199,8)),
			8508 => std_logic_vector(to_unsigned( 247,8)),
			8509 => std_logic_vector(to_unsigned( 122,8)),
			8510 => std_logic_vector(to_unsigned( 67,8)),
			8511 => std_logic_vector(to_unsigned( 211,8)),
			8512 => std_logic_vector(to_unsigned( 123,8)),
			8513 => std_logic_vector(to_unsigned( 119,8)),
			8514 => std_logic_vector(to_unsigned( 73,8)),
			8515 => std_logic_vector(to_unsigned( 134,8)),
			8516 => std_logic_vector(to_unsigned( 169,8)),
			8517 => std_logic_vector(to_unsigned( 34,8)),
			8518 => std_logic_vector(to_unsigned( 129,8)),
			8519 => std_logic_vector(to_unsigned( 113,8)),
			8520 => std_logic_vector(to_unsigned( 192,8)),
			8521 => std_logic_vector(to_unsigned( 173,8)),
			8522 => std_logic_vector(to_unsigned( 170,8)),
			8523 => std_logic_vector(to_unsigned( 170,8)),
			8524 => std_logic_vector(to_unsigned( 5,8)),
			8525 => std_logic_vector(to_unsigned( 167,8)),
			8526 => std_logic_vector(to_unsigned( 160,8)),
			8527 => std_logic_vector(to_unsigned( 231,8)),
			8528 => std_logic_vector(to_unsigned( 198,8)),
			8529 => std_logic_vector(to_unsigned( 71,8)),
			8530 => std_logic_vector(to_unsigned( 44,8)),
			8531 => std_logic_vector(to_unsigned( 152,8)),
			8532 => std_logic_vector(to_unsigned( 244,8)),
			8533 => std_logic_vector(to_unsigned( 252,8)),
			8534 => std_logic_vector(to_unsigned( 194,8)),
			8535 => std_logic_vector(to_unsigned( 174,8)),
			8536 => std_logic_vector(to_unsigned( 105,8)),
			8537 => std_logic_vector(to_unsigned( 172,8)),
			8538 => std_logic_vector(to_unsigned( 112,8)),
			8539 => std_logic_vector(to_unsigned( 155,8)),
			8540 => std_logic_vector(to_unsigned( 26,8)),
			8541 => std_logic_vector(to_unsigned( 117,8)),
			8542 => std_logic_vector(to_unsigned( 174,8)),
			8543 => std_logic_vector(to_unsigned( 184,8)),
			8544 => std_logic_vector(to_unsigned( 60,8)),
			8545 => std_logic_vector(to_unsigned( 79,8)),
			8546 => std_logic_vector(to_unsigned( 231,8)),
			8547 => std_logic_vector(to_unsigned( 17,8)),
			8548 => std_logic_vector(to_unsigned( 129,8)),
			8549 => std_logic_vector(to_unsigned( 34,8)),
			8550 => std_logic_vector(to_unsigned( 165,8)),
			8551 => std_logic_vector(to_unsigned( 152,8)),
			8552 => std_logic_vector(to_unsigned( 154,8)),
			8553 => std_logic_vector(to_unsigned( 236,8)),
			8554 => std_logic_vector(to_unsigned( 106,8)),
			8555 => std_logic_vector(to_unsigned( 6,8)),
			8556 => std_logic_vector(to_unsigned( 233,8)),
			8557 => std_logic_vector(to_unsigned( 104,8)),
			8558 => std_logic_vector(to_unsigned( 89,8)),
			8559 => std_logic_vector(to_unsigned( 61,8)),
			8560 => std_logic_vector(to_unsigned( 59,8)),
			8561 => std_logic_vector(to_unsigned( 177,8)),
			8562 => std_logic_vector(to_unsigned( 189,8)),
			8563 => std_logic_vector(to_unsigned( 126,8)),
			8564 => std_logic_vector(to_unsigned( 221,8)),
			8565 => std_logic_vector(to_unsigned( 178,8)),
			8566 => std_logic_vector(to_unsigned( 93,8)),
			8567 => std_logic_vector(to_unsigned( 211,8)),
			8568 => std_logic_vector(to_unsigned( 189,8)),
			8569 => std_logic_vector(to_unsigned( 101,8)),
			8570 => std_logic_vector(to_unsigned( 42,8)),
			8571 => std_logic_vector(to_unsigned( 142,8)),
			8572 => std_logic_vector(to_unsigned( 51,8)),
			8573 => std_logic_vector(to_unsigned( 167,8)),
			8574 => std_logic_vector(to_unsigned( 233,8)),
			8575 => std_logic_vector(to_unsigned( 134,8)),
			8576 => std_logic_vector(to_unsigned( 223,8)),
			8577 => std_logic_vector(to_unsigned( 158,8)),
			8578 => std_logic_vector(to_unsigned( 249,8)),
			8579 => std_logic_vector(to_unsigned( 108,8)),
			8580 => std_logic_vector(to_unsigned( 133,8)),
			8581 => std_logic_vector(to_unsigned( 151,8)),
			8582 => std_logic_vector(to_unsigned( 85,8)),
			8583 => std_logic_vector(to_unsigned( 252,8)),
			8584 => std_logic_vector(to_unsigned( 77,8)),
			8585 => std_logic_vector(to_unsigned( 165,8)),
			8586 => std_logic_vector(to_unsigned( 23,8)),
			8587 => std_logic_vector(to_unsigned( 242,8)),
			8588 => std_logic_vector(to_unsigned( 188,8)),
			8589 => std_logic_vector(to_unsigned( 248,8)),
			8590 => std_logic_vector(to_unsigned( 174,8)),
			8591 => std_logic_vector(to_unsigned( 178,8)),
			8592 => std_logic_vector(to_unsigned( 92,8)),
			8593 => std_logic_vector(to_unsigned( 157,8)),
			8594 => std_logic_vector(to_unsigned( 30,8)),
			8595 => std_logic_vector(to_unsigned( 203,8)),
			8596 => std_logic_vector(to_unsigned( 87,8)),
			8597 => std_logic_vector(to_unsigned( 144,8)),
			8598 => std_logic_vector(to_unsigned( 93,8)),
			8599 => std_logic_vector(to_unsigned( 14,8)),
			8600 => std_logic_vector(to_unsigned( 255,8)),
			8601 => std_logic_vector(to_unsigned( 31,8)),
			8602 => std_logic_vector(to_unsigned( 73,8)),
			8603 => std_logic_vector(to_unsigned( 93,8)),
			8604 => std_logic_vector(to_unsigned( 187,8)),
			8605 => std_logic_vector(to_unsigned( 161,8)),
			8606 => std_logic_vector(to_unsigned( 13,8)),
			8607 => std_logic_vector(to_unsigned( 223,8)),
			8608 => std_logic_vector(to_unsigned( 118,8)),
			8609 => std_logic_vector(to_unsigned( 75,8)),
			8610 => std_logic_vector(to_unsigned( 30,8)),
			8611 => std_logic_vector(to_unsigned( 229,8)),
			8612 => std_logic_vector(to_unsigned( 88,8)),
			8613 => std_logic_vector(to_unsigned( 128,8)),
			8614 => std_logic_vector(to_unsigned( 194,8)),
			8615 => std_logic_vector(to_unsigned( 53,8)),
			8616 => std_logic_vector(to_unsigned( 129,8)),
			8617 => std_logic_vector(to_unsigned( 161,8)),
			8618 => std_logic_vector(to_unsigned( 147,8)),
			8619 => std_logic_vector(to_unsigned( 50,8)),
			8620 => std_logic_vector(to_unsigned( 168,8)),
			8621 => std_logic_vector(to_unsigned( 249,8)),
			8622 => std_logic_vector(to_unsigned( 18,8)),
			8623 => std_logic_vector(to_unsigned( 116,8)),
			8624 => std_logic_vector(to_unsigned( 4,8)),
			8625 => std_logic_vector(to_unsigned( 105,8)),
			8626 => std_logic_vector(to_unsigned( 29,8)),
			8627 => std_logic_vector(to_unsigned( 105,8)),
			8628 => std_logic_vector(to_unsigned( 73,8)),
			8629 => std_logic_vector(to_unsigned( 198,8)),
			8630 => std_logic_vector(to_unsigned( 174,8)),
			8631 => std_logic_vector(to_unsigned( 192,8)),
			8632 => std_logic_vector(to_unsigned( 48,8)),
			8633 => std_logic_vector(to_unsigned( 114,8)),
			8634 => std_logic_vector(to_unsigned( 20,8)),
			8635 => std_logic_vector(to_unsigned( 40,8)),
			8636 => std_logic_vector(to_unsigned( 251,8)),
			8637 => std_logic_vector(to_unsigned( 206,8)),
			8638 => std_logic_vector(to_unsigned( 119,8)),
			8639 => std_logic_vector(to_unsigned( 187,8)),
			8640 => std_logic_vector(to_unsigned( 165,8)),
			8641 => std_logic_vector(to_unsigned( 246,8)),
			8642 => std_logic_vector(to_unsigned( 240,8)),
			8643 => std_logic_vector(to_unsigned( 54,8)),
			8644 => std_logic_vector(to_unsigned( 162,8)),
			8645 => std_logic_vector(to_unsigned( 245,8)),
			8646 => std_logic_vector(to_unsigned( 5,8)),
			8647 => std_logic_vector(to_unsigned( 75,8)),
			8648 => std_logic_vector(to_unsigned( 255,8)),
			8649 => std_logic_vector(to_unsigned( 130,8)),
			8650 => std_logic_vector(to_unsigned( 10,8)),
			8651 => std_logic_vector(to_unsigned( 117,8)),
			8652 => std_logic_vector(to_unsigned( 174,8)),
			8653 => std_logic_vector(to_unsigned( 156,8)),
			8654 => std_logic_vector(to_unsigned( 215,8)),
			8655 => std_logic_vector(to_unsigned( 76,8)),
			8656 => std_logic_vector(to_unsigned( 120,8)),
			8657 => std_logic_vector(to_unsigned( 51,8)),
			8658 => std_logic_vector(to_unsigned( 128,8)),
			8659 => std_logic_vector(to_unsigned( 20,8)),
			8660 => std_logic_vector(to_unsigned( 243,8)),
			8661 => std_logic_vector(to_unsigned( 84,8)),
			8662 => std_logic_vector(to_unsigned( 200,8)),
			8663 => std_logic_vector(to_unsigned( 1,8)),
			8664 => std_logic_vector(to_unsigned( 242,8)),
			8665 => std_logic_vector(to_unsigned( 116,8)),
			8666 => std_logic_vector(to_unsigned( 127,8)),
			8667 => std_logic_vector(to_unsigned( 236,8)),
			8668 => std_logic_vector(to_unsigned( 81,8)),
			8669 => std_logic_vector(to_unsigned( 185,8)),
			8670 => std_logic_vector(to_unsigned( 81,8)),
			8671 => std_logic_vector(to_unsigned( 113,8)),
			8672 => std_logic_vector(to_unsigned( 229,8)),
			8673 => std_logic_vector(to_unsigned( 222,8)),
			8674 => std_logic_vector(to_unsigned( 84,8)),
			8675 => std_logic_vector(to_unsigned( 232,8)),
			8676 => std_logic_vector(to_unsigned( 99,8)),
			8677 => std_logic_vector(to_unsigned( 222,8)),
			8678 => std_logic_vector(to_unsigned( 123,8)),
			8679 => std_logic_vector(to_unsigned( 195,8)),
			8680 => std_logic_vector(to_unsigned( 187,8)),
			8681 => std_logic_vector(to_unsigned( 196,8)),
			8682 => std_logic_vector(to_unsigned( 175,8)),
			8683 => std_logic_vector(to_unsigned( 172,8)),
			8684 => std_logic_vector(to_unsigned( 236,8)),
			8685 => std_logic_vector(to_unsigned( 211,8)),
			8686 => std_logic_vector(to_unsigned( 60,8)),
			8687 => std_logic_vector(to_unsigned( 108,8)),
			8688 => std_logic_vector(to_unsigned( 100,8)),
			8689 => std_logic_vector(to_unsigned( 165,8)),
			8690 => std_logic_vector(to_unsigned( 158,8)),
			8691 => std_logic_vector(to_unsigned( 134,8)),
			8692 => std_logic_vector(to_unsigned( 117,8)),
			8693 => std_logic_vector(to_unsigned( 114,8)),
			8694 => std_logic_vector(to_unsigned( 150,8)),
			8695 => std_logic_vector(to_unsigned( 224,8)),
			8696 => std_logic_vector(to_unsigned( 162,8)),
			8697 => std_logic_vector(to_unsigned( 76,8)),
			8698 => std_logic_vector(to_unsigned( 114,8)),
			8699 => std_logic_vector(to_unsigned( 91,8)),
			8700 => std_logic_vector(to_unsigned( 238,8)),
			8701 => std_logic_vector(to_unsigned( 140,8)),
			8702 => std_logic_vector(to_unsigned( 209,8)),
			8703 => std_logic_vector(to_unsigned( 28,8)),
			8704 => std_logic_vector(to_unsigned( 52,8)),
			8705 => std_logic_vector(to_unsigned( 102,8)),
			8706 => std_logic_vector(to_unsigned( 104,8)),
			8707 => std_logic_vector(to_unsigned( 22,8)),
			8708 => std_logic_vector(to_unsigned( 14,8)),
			8709 => std_logic_vector(to_unsigned( 51,8)),
			8710 => std_logic_vector(to_unsigned( 237,8)),
			8711 => std_logic_vector(to_unsigned( 14,8)),
			8712 => std_logic_vector(to_unsigned( 2,8)),
			8713 => std_logic_vector(to_unsigned( 193,8)),
			8714 => std_logic_vector(to_unsigned( 246,8)),
			8715 => std_logic_vector(to_unsigned( 131,8)),
			8716 => std_logic_vector(to_unsigned( 111,8)),
			8717 => std_logic_vector(to_unsigned( 108,8)),
			8718 => std_logic_vector(to_unsigned( 228,8)),
			8719 => std_logic_vector(to_unsigned( 34,8)),
			8720 => std_logic_vector(to_unsigned( 2,8)),
			8721 => std_logic_vector(to_unsigned( 54,8)),
			8722 => std_logic_vector(to_unsigned( 172,8)),
			8723 => std_logic_vector(to_unsigned( 36,8)),
			8724 => std_logic_vector(to_unsigned( 113,8)),
			8725 => std_logic_vector(to_unsigned( 43,8)),
			8726 => std_logic_vector(to_unsigned( 215,8)),
			8727 => std_logic_vector(to_unsigned( 132,8)),
			8728 => std_logic_vector(to_unsigned( 0,8)),
			8729 => std_logic_vector(to_unsigned( 206,8)),
			8730 => std_logic_vector(to_unsigned( 165,8)),
			8731 => std_logic_vector(to_unsigned( 75,8)),
			8732 => std_logic_vector(to_unsigned( 92,8)),
			8733 => std_logic_vector(to_unsigned( 70,8)),
			8734 => std_logic_vector(to_unsigned( 7,8)),
			8735 => std_logic_vector(to_unsigned( 226,8)),
			8736 => std_logic_vector(to_unsigned( 36,8)),
			8737 => std_logic_vector(to_unsigned( 218,8)),
			8738 => std_logic_vector(to_unsigned( 105,8)),
			8739 => std_logic_vector(to_unsigned( 81,8)),
			8740 => std_logic_vector(to_unsigned( 247,8)),
			8741 => std_logic_vector(to_unsigned( 25,8)),
			8742 => std_logic_vector(to_unsigned( 78,8)),
			8743 => std_logic_vector(to_unsigned( 107,8)),
			8744 => std_logic_vector(to_unsigned( 105,8)),
			8745 => std_logic_vector(to_unsigned( 203,8)),
			8746 => std_logic_vector(to_unsigned( 58,8)),
			8747 => std_logic_vector(to_unsigned( 6,8)),
			8748 => std_logic_vector(to_unsigned( 101,8)),
			8749 => std_logic_vector(to_unsigned( 223,8)),
			8750 => std_logic_vector(to_unsigned( 37,8)),
			8751 => std_logic_vector(to_unsigned( 227,8)),
			8752 => std_logic_vector(to_unsigned( 163,8)),
			8753 => std_logic_vector(to_unsigned( 52,8)),
			8754 => std_logic_vector(to_unsigned( 120,8)),
			8755 => std_logic_vector(to_unsigned( 78,8)),
			8756 => std_logic_vector(to_unsigned( 165,8)),
			8757 => std_logic_vector(to_unsigned( 40,8)),
			8758 => std_logic_vector(to_unsigned( 187,8)),
			8759 => std_logic_vector(to_unsigned( 246,8)),
			8760 => std_logic_vector(to_unsigned( 225,8)),
			8761 => std_logic_vector(to_unsigned( 156,8)),
			8762 => std_logic_vector(to_unsigned( 92,8)),
			8763 => std_logic_vector(to_unsigned( 4,8)),
			8764 => std_logic_vector(to_unsigned( 252,8)),
			8765 => std_logic_vector(to_unsigned( 89,8)),
			8766 => std_logic_vector(to_unsigned( 43,8)),
			8767 => std_logic_vector(to_unsigned( 254,8)),
			8768 => std_logic_vector(to_unsigned( 155,8)),
			8769 => std_logic_vector(to_unsigned( 39,8)),
			8770 => std_logic_vector(to_unsigned( 58,8)),
			8771 => std_logic_vector(to_unsigned( 134,8)),
			8772 => std_logic_vector(to_unsigned( 91,8)),
			8773 => std_logic_vector(to_unsigned( 250,8)),
			8774 => std_logic_vector(to_unsigned( 249,8)),
			8775 => std_logic_vector(to_unsigned( 32,8)),
			8776 => std_logic_vector(to_unsigned( 194,8)),
			8777 => std_logic_vector(to_unsigned( 185,8)),
			8778 => std_logic_vector(to_unsigned( 238,8)),
			8779 => std_logic_vector(to_unsigned( 108,8)),
			8780 => std_logic_vector(to_unsigned( 22,8)),
			8781 => std_logic_vector(to_unsigned( 94,8)),
			8782 => std_logic_vector(to_unsigned( 229,8)),
			8783 => std_logic_vector(to_unsigned( 13,8)),
			8784 => std_logic_vector(to_unsigned( 33,8)),
			8785 => std_logic_vector(to_unsigned( 29,8)),
			8786 => std_logic_vector(to_unsigned( 81,8)),
			8787 => std_logic_vector(to_unsigned( 14,8)),
			8788 => std_logic_vector(to_unsigned( 207,8)),
			8789 => std_logic_vector(to_unsigned( 104,8)),
			8790 => std_logic_vector(to_unsigned( 167,8)),
			8791 => std_logic_vector(to_unsigned( 45,8)),
			8792 => std_logic_vector(to_unsigned( 138,8)),
			8793 => std_logic_vector(to_unsigned( 139,8)),
			8794 => std_logic_vector(to_unsigned( 169,8)),
			8795 => std_logic_vector(to_unsigned( 38,8)),
			8796 => std_logic_vector(to_unsigned( 71,8)),
			8797 => std_logic_vector(to_unsigned( 153,8)),
			8798 => std_logic_vector(to_unsigned( 96,8)),
			8799 => std_logic_vector(to_unsigned( 98,8)),
			8800 => std_logic_vector(to_unsigned( 200,8)),
			8801 => std_logic_vector(to_unsigned( 172,8)),
			8802 => std_logic_vector(to_unsigned( 170,8)),
			8803 => std_logic_vector(to_unsigned( 125,8)),
			8804 => std_logic_vector(to_unsigned( 58,8)),
			8805 => std_logic_vector(to_unsigned( 242,8)),
			8806 => std_logic_vector(to_unsigned( 40,8)),
			8807 => std_logic_vector(to_unsigned( 84,8)),
			8808 => std_logic_vector(to_unsigned( 26,8)),
			8809 => std_logic_vector(to_unsigned( 210,8)),
			8810 => std_logic_vector(to_unsigned( 226,8)),
			8811 => std_logic_vector(to_unsigned( 131,8)),
			8812 => std_logic_vector(to_unsigned( 166,8)),
			8813 => std_logic_vector(to_unsigned( 118,8)),
			8814 => std_logic_vector(to_unsigned( 14,8)),
			8815 => std_logic_vector(to_unsigned( 52,8)),
			8816 => std_logic_vector(to_unsigned( 223,8)),
			8817 => std_logic_vector(to_unsigned( 244,8)),
			8818 => std_logic_vector(to_unsigned( 195,8)),
			8819 => std_logic_vector(to_unsigned( 57,8)),
			8820 => std_logic_vector(to_unsigned( 101,8)),
			8821 => std_logic_vector(to_unsigned( 31,8)),
			8822 => std_logic_vector(to_unsigned( 160,8)),
			8823 => std_logic_vector(to_unsigned( 45,8)),
			8824 => std_logic_vector(to_unsigned( 140,8)),
			8825 => std_logic_vector(to_unsigned( 29,8)),
			8826 => std_logic_vector(to_unsigned( 139,8)),
			8827 => std_logic_vector(to_unsigned( 8,8)),
			8828 => std_logic_vector(to_unsigned( 28,8)),
			8829 => std_logic_vector(to_unsigned( 158,8)),
			8830 => std_logic_vector(to_unsigned( 184,8)),
			8831 => std_logic_vector(to_unsigned( 127,8)),
			8832 => std_logic_vector(to_unsigned( 113,8)),
			8833 => std_logic_vector(to_unsigned( 62,8)),
			8834 => std_logic_vector(to_unsigned( 12,8)),
			8835 => std_logic_vector(to_unsigned( 181,8)),
			8836 => std_logic_vector(to_unsigned( 24,8)),
			8837 => std_logic_vector(to_unsigned( 140,8)),
			8838 => std_logic_vector(to_unsigned( 168,8)),
			8839 => std_logic_vector(to_unsigned( 62,8)),
			8840 => std_logic_vector(to_unsigned( 53,8)),
			8841 => std_logic_vector(to_unsigned( 219,8)),
			8842 => std_logic_vector(to_unsigned( 158,8)),
			8843 => std_logic_vector(to_unsigned( 142,8)),
			8844 => std_logic_vector(to_unsigned( 140,8)),
			8845 => std_logic_vector(to_unsigned( 27,8)),
			8846 => std_logic_vector(to_unsigned( 218,8)),
			8847 => std_logic_vector(to_unsigned( 5,8)),
			8848 => std_logic_vector(to_unsigned( 148,8)),
			8849 => std_logic_vector(to_unsigned( 236,8)),
			8850 => std_logic_vector(to_unsigned( 100,8)),
			8851 => std_logic_vector(to_unsigned( 9,8)),
			8852 => std_logic_vector(to_unsigned( 149,8)),
			8853 => std_logic_vector(to_unsigned( 174,8)),
			8854 => std_logic_vector(to_unsigned( 13,8)),
			8855 => std_logic_vector(to_unsigned( 152,8)),
			8856 => std_logic_vector(to_unsigned( 10,8)),
			8857 => std_logic_vector(to_unsigned( 59,8)),
			8858 => std_logic_vector(to_unsigned( 85,8)),
			8859 => std_logic_vector(to_unsigned( 109,8)),
			8860 => std_logic_vector(to_unsigned( 207,8)),
			8861 => std_logic_vector(to_unsigned( 124,8)),
			8862 => std_logic_vector(to_unsigned( 147,8)),
			8863 => std_logic_vector(to_unsigned( 218,8)),
			8864 => std_logic_vector(to_unsigned( 175,8)),
			8865 => std_logic_vector(to_unsigned( 186,8)),
			8866 => std_logic_vector(to_unsigned( 127,8)),
			8867 => std_logic_vector(to_unsigned( 5,8)),
			8868 => std_logic_vector(to_unsigned( 248,8)),
			8869 => std_logic_vector(to_unsigned( 37,8)),
			8870 => std_logic_vector(to_unsigned( 153,8)),
			8871 => std_logic_vector(to_unsigned( 40,8)),
			8872 => std_logic_vector(to_unsigned( 193,8)),
			8873 => std_logic_vector(to_unsigned( 166,8)),
			8874 => std_logic_vector(to_unsigned( 204,8)),
			8875 => std_logic_vector(to_unsigned( 128,8)),
			8876 => std_logic_vector(to_unsigned( 46,8)),
			8877 => std_logic_vector(to_unsigned( 31,8)),
			8878 => std_logic_vector(to_unsigned( 44,8)),
			8879 => std_logic_vector(to_unsigned( 83,8)),
			8880 => std_logic_vector(to_unsigned( 11,8)),
			8881 => std_logic_vector(to_unsigned( 68,8)),
			8882 => std_logic_vector(to_unsigned( 99,8)),
			8883 => std_logic_vector(to_unsigned( 40,8)),
			8884 => std_logic_vector(to_unsigned( 127,8)),
			8885 => std_logic_vector(to_unsigned( 29,8)),
			8886 => std_logic_vector(to_unsigned( 101,8)),
			8887 => std_logic_vector(to_unsigned( 50,8)),
			8888 => std_logic_vector(to_unsigned( 253,8)),
			8889 => std_logic_vector(to_unsigned( 103,8)),
			8890 => std_logic_vector(to_unsigned( 236,8)),
			8891 => std_logic_vector(to_unsigned( 65,8)),
			8892 => std_logic_vector(to_unsigned( 60,8)),
			8893 => std_logic_vector(to_unsigned( 49,8)),
			8894 => std_logic_vector(to_unsigned( 152,8)),
			8895 => std_logic_vector(to_unsigned( 204,8)),
			8896 => std_logic_vector(to_unsigned( 146,8)),
			8897 => std_logic_vector(to_unsigned( 94,8)),
			8898 => std_logic_vector(to_unsigned( 147,8)),
			8899 => std_logic_vector(to_unsigned( 58,8)),
			8900 => std_logic_vector(to_unsigned( 48,8)),
			8901 => std_logic_vector(to_unsigned( 33,8)),
			8902 => std_logic_vector(to_unsigned( 38,8)),
			8903 => std_logic_vector(to_unsigned( 147,8)),
			8904 => std_logic_vector(to_unsigned( 111,8)),
			8905 => std_logic_vector(to_unsigned( 217,8)),
			8906 => std_logic_vector(to_unsigned( 107,8)),
			8907 => std_logic_vector(to_unsigned( 17,8)),
			8908 => std_logic_vector(to_unsigned( 220,8)),
			8909 => std_logic_vector(to_unsigned( 40,8)),
			8910 => std_logic_vector(to_unsigned( 243,8)),
			8911 => std_logic_vector(to_unsigned( 2,8)),
			8912 => std_logic_vector(to_unsigned( 179,8)),
			8913 => std_logic_vector(to_unsigned( 11,8)),
			8914 => std_logic_vector(to_unsigned( 7,8)),
			8915 => std_logic_vector(to_unsigned( 91,8)),
			8916 => std_logic_vector(to_unsigned( 45,8)),
			8917 => std_logic_vector(to_unsigned( 154,8)),
			8918 => std_logic_vector(to_unsigned( 76,8)),
			8919 => std_logic_vector(to_unsigned( 171,8)),
			8920 => std_logic_vector(to_unsigned( 231,8)),
			8921 => std_logic_vector(to_unsigned( 196,8)),
			8922 => std_logic_vector(to_unsigned( 131,8)),
			8923 => std_logic_vector(to_unsigned( 110,8)),
			8924 => std_logic_vector(to_unsigned( 216,8)),
			8925 => std_logic_vector(to_unsigned( 134,8)),
			8926 => std_logic_vector(to_unsigned( 33,8)),
			8927 => std_logic_vector(to_unsigned( 2,8)),
			8928 => std_logic_vector(to_unsigned( 192,8)),
			8929 => std_logic_vector(to_unsigned( 144,8)),
			8930 => std_logic_vector(to_unsigned( 204,8)),
			8931 => std_logic_vector(to_unsigned( 221,8)),
			8932 => std_logic_vector(to_unsigned( 18,8)),
			8933 => std_logic_vector(to_unsigned( 233,8)),
			8934 => std_logic_vector(to_unsigned( 200,8)),
			8935 => std_logic_vector(to_unsigned( 193,8)),
			8936 => std_logic_vector(to_unsigned( 6,8)),
			8937 => std_logic_vector(to_unsigned( 75,8)),
			8938 => std_logic_vector(to_unsigned( 121,8)),
			8939 => std_logic_vector(to_unsigned( 216,8)),
			8940 => std_logic_vector(to_unsigned( 188,8)),
			8941 => std_logic_vector(to_unsigned( 136,8)),
			8942 => std_logic_vector(to_unsigned( 30,8)),
			8943 => std_logic_vector(to_unsigned( 127,8)),
			8944 => std_logic_vector(to_unsigned( 51,8)),
			8945 => std_logic_vector(to_unsigned( 255,8)),
			8946 => std_logic_vector(to_unsigned( 195,8)),
			8947 => std_logic_vector(to_unsigned( 235,8)),
			8948 => std_logic_vector(to_unsigned( 121,8)),
			8949 => std_logic_vector(to_unsigned( 128,8)),
			8950 => std_logic_vector(to_unsigned( 205,8)),
			8951 => std_logic_vector(to_unsigned( 45,8)),
			8952 => std_logic_vector(to_unsigned( 220,8)),
			8953 => std_logic_vector(to_unsigned( 190,8)),
			8954 => std_logic_vector(to_unsigned( 195,8)),
			8955 => std_logic_vector(to_unsigned( 190,8)),
			8956 => std_logic_vector(to_unsigned( 240,8)),
			8957 => std_logic_vector(to_unsigned( 124,8)),
			8958 => std_logic_vector(to_unsigned( 66,8)),
			8959 => std_logic_vector(to_unsigned( 46,8)),
			8960 => std_logic_vector(to_unsigned( 198,8)),
			8961 => std_logic_vector(to_unsigned( 148,8)),
			8962 => std_logic_vector(to_unsigned( 252,8)),
			8963 => std_logic_vector(to_unsigned( 75,8)),
			8964 => std_logic_vector(to_unsigned( 23,8)),
			8965 => std_logic_vector(to_unsigned( 30,8)),
			8966 => std_logic_vector(to_unsigned( 37,8)),
			8967 => std_logic_vector(to_unsigned( 2,8)),
			8968 => std_logic_vector(to_unsigned( 189,8)),
			8969 => std_logic_vector(to_unsigned( 73,8)),
			8970 => std_logic_vector(to_unsigned( 116,8)),
			8971 => std_logic_vector(to_unsigned( 246,8)),
			8972 => std_logic_vector(to_unsigned( 48,8)),
			8973 => std_logic_vector(to_unsigned( 122,8)),
			8974 => std_logic_vector(to_unsigned( 61,8)),
			8975 => std_logic_vector(to_unsigned( 177,8)),
			8976 => std_logic_vector(to_unsigned( 73,8)),
			8977 => std_logic_vector(to_unsigned( 125,8)),
			8978 => std_logic_vector(to_unsigned( 126,8)),
			8979 => std_logic_vector(to_unsigned( 247,8)),
			8980 => std_logic_vector(to_unsigned( 122,8)),
			8981 => std_logic_vector(to_unsigned( 81,8)),
			8982 => std_logic_vector(to_unsigned( 65,8)),
			8983 => std_logic_vector(to_unsigned( 226,8)),
			8984 => std_logic_vector(to_unsigned( 138,8)),
			8985 => std_logic_vector(to_unsigned( 25,8)),
			8986 => std_logic_vector(to_unsigned( 242,8)),
			8987 => std_logic_vector(to_unsigned( 23,8)),
			8988 => std_logic_vector(to_unsigned( 231,8)),
			8989 => std_logic_vector(to_unsigned( 148,8)),
			8990 => std_logic_vector(to_unsigned( 25,8)),
			8991 => std_logic_vector(to_unsigned( 203,8)),
			8992 => std_logic_vector(to_unsigned( 216,8)),
			8993 => std_logic_vector(to_unsigned( 130,8)),
			8994 => std_logic_vector(to_unsigned( 135,8)),
			8995 => std_logic_vector(to_unsigned( 63,8)),
			8996 => std_logic_vector(to_unsigned( 216,8)),
			8997 => std_logic_vector(to_unsigned( 201,8)),
			8998 => std_logic_vector(to_unsigned( 36,8)),
			8999 => std_logic_vector(to_unsigned( 251,8)),
			9000 => std_logic_vector(to_unsigned( 196,8)),
			9001 => std_logic_vector(to_unsigned( 192,8)),
			9002 => std_logic_vector(to_unsigned( 217,8)),
			9003 => std_logic_vector(to_unsigned( 190,8)),
			9004 => std_logic_vector(to_unsigned( 153,8)),
			9005 => std_logic_vector(to_unsigned( 51,8)),
			9006 => std_logic_vector(to_unsigned( 129,8)),
			9007 => std_logic_vector(to_unsigned( 246,8)),
			9008 => std_logic_vector(to_unsigned( 130,8)),
			9009 => std_logic_vector(to_unsigned( 94,8)),
			9010 => std_logic_vector(to_unsigned( 82,8)),
			9011 => std_logic_vector(to_unsigned( 19,8)),
			9012 => std_logic_vector(to_unsigned( 59,8)),
			9013 => std_logic_vector(to_unsigned( 46,8)),
			9014 => std_logic_vector(to_unsigned( 188,8)),
			9015 => std_logic_vector(to_unsigned( 48,8)),
			9016 => std_logic_vector(to_unsigned( 6,8)),
			9017 => std_logic_vector(to_unsigned( 141,8)),
			9018 => std_logic_vector(to_unsigned( 53,8)),
			9019 => std_logic_vector(to_unsigned( 189,8)),
			9020 => std_logic_vector(to_unsigned( 216,8)),
			9021 => std_logic_vector(to_unsigned( 237,8)),
			9022 => std_logic_vector(to_unsigned( 2,8)),
			9023 => std_logic_vector(to_unsigned( 115,8)),
			9024 => std_logic_vector(to_unsigned( 39,8)),
			9025 => std_logic_vector(to_unsigned( 54,8)),
			9026 => std_logic_vector(to_unsigned( 189,8)),
			9027 => std_logic_vector(to_unsigned( 147,8)),
			9028 => std_logic_vector(to_unsigned( 41,8)),
			9029 => std_logic_vector(to_unsigned( 165,8)),
			9030 => std_logic_vector(to_unsigned( 26,8)),
			9031 => std_logic_vector(to_unsigned( 72,8)),
			9032 => std_logic_vector(to_unsigned( 85,8)),
			9033 => std_logic_vector(to_unsigned( 115,8)),
			9034 => std_logic_vector(to_unsigned( 237,8)),
			9035 => std_logic_vector(to_unsigned( 238,8)),
			9036 => std_logic_vector(to_unsigned( 189,8)),
			9037 => std_logic_vector(to_unsigned( 8,8)),
			9038 => std_logic_vector(to_unsigned( 179,8)),
			9039 => std_logic_vector(to_unsigned( 6,8)),
			9040 => std_logic_vector(to_unsigned( 59,8)),
			9041 => std_logic_vector(to_unsigned( 166,8)),
			9042 => std_logic_vector(to_unsigned( 121,8)),
			9043 => std_logic_vector(to_unsigned( 43,8)),
			9044 => std_logic_vector(to_unsigned( 217,8)),
			9045 => std_logic_vector(to_unsigned( 134,8)),
			9046 => std_logic_vector(to_unsigned( 131,8)),
			9047 => std_logic_vector(to_unsigned( 165,8)),
			9048 => std_logic_vector(to_unsigned( 240,8)),
			9049 => std_logic_vector(to_unsigned( 11,8)),
			9050 => std_logic_vector(to_unsigned( 32,8)),
			9051 => std_logic_vector(to_unsigned( 43,8)),
			9052 => std_logic_vector(to_unsigned( 179,8)),
			9053 => std_logic_vector(to_unsigned( 166,8)),
			9054 => std_logic_vector(to_unsigned( 112,8)),
			9055 => std_logic_vector(to_unsigned( 64,8)),
			9056 => std_logic_vector(to_unsigned( 113,8)),
			9057 => std_logic_vector(to_unsigned( 193,8)),
			9058 => std_logic_vector(to_unsigned( 39,8)),
			9059 => std_logic_vector(to_unsigned( 81,8)),
			9060 => std_logic_vector(to_unsigned( 103,8)),
			9061 => std_logic_vector(to_unsigned( 43,8)),
			9062 => std_logic_vector(to_unsigned( 223,8)),
			9063 => std_logic_vector(to_unsigned( 191,8)),
			9064 => std_logic_vector(to_unsigned( 82,8)),
			9065 => std_logic_vector(to_unsigned( 26,8)),
			9066 => std_logic_vector(to_unsigned( 52,8)),
			9067 => std_logic_vector(to_unsigned( 56,8)),
			9068 => std_logic_vector(to_unsigned( 209,8)),
			9069 => std_logic_vector(to_unsigned( 203,8)),
			9070 => std_logic_vector(to_unsigned( 12,8)),
			9071 => std_logic_vector(to_unsigned( 17,8)),
			9072 => std_logic_vector(to_unsigned( 141,8)),
			9073 => std_logic_vector(to_unsigned( 180,8)),
			9074 => std_logic_vector(to_unsigned( 152,8)),
			9075 => std_logic_vector(to_unsigned( 105,8)),
			9076 => std_logic_vector(to_unsigned( 179,8)),
			9077 => std_logic_vector(to_unsigned( 132,8)),
			9078 => std_logic_vector(to_unsigned( 181,8)),
			9079 => std_logic_vector(to_unsigned( 167,8)),
			9080 => std_logic_vector(to_unsigned( 70,8)),
			9081 => std_logic_vector(to_unsigned( 67,8)),
			9082 => std_logic_vector(to_unsigned( 52,8)),
			9083 => std_logic_vector(to_unsigned( 160,8)),
			9084 => std_logic_vector(to_unsigned( 209,8)),
			9085 => std_logic_vector(to_unsigned( 250,8)),
			9086 => std_logic_vector(to_unsigned( 167,8)),
			9087 => std_logic_vector(to_unsigned( 93,8)),
			9088 => std_logic_vector(to_unsigned( 23,8)),
			9089 => std_logic_vector(to_unsigned( 76,8)),
			9090 => std_logic_vector(to_unsigned( 37,8)),
			9091 => std_logic_vector(to_unsigned( 164,8)),
			9092 => std_logic_vector(to_unsigned( 130,8)),
			9093 => std_logic_vector(to_unsigned( 83,8)),
			9094 => std_logic_vector(to_unsigned( 121,8)),
			9095 => std_logic_vector(to_unsigned( 46,8)),
			9096 => std_logic_vector(to_unsigned( 35,8)),
			9097 => std_logic_vector(to_unsigned( 172,8)),
			9098 => std_logic_vector(to_unsigned( 207,8)),
			9099 => std_logic_vector(to_unsigned( 15,8)),
			9100 => std_logic_vector(to_unsigned( 4,8)),
			9101 => std_logic_vector(to_unsigned( 151,8)),
			9102 => std_logic_vector(to_unsigned( 238,8)),
			9103 => std_logic_vector(to_unsigned( 130,8)),
			9104 => std_logic_vector(to_unsigned( 91,8)),
			9105 => std_logic_vector(to_unsigned( 206,8)),
			9106 => std_logic_vector(to_unsigned( 112,8)),
			9107 => std_logic_vector(to_unsigned( 119,8)),
			9108 => std_logic_vector(to_unsigned( 140,8)),
			9109 => std_logic_vector(to_unsigned( 30,8)),
			9110 => std_logic_vector(to_unsigned( 1,8)),
			9111 => std_logic_vector(to_unsigned( 222,8)),
			9112 => std_logic_vector(to_unsigned( 248,8)),
			9113 => std_logic_vector(to_unsigned( 211,8)),
			9114 => std_logic_vector(to_unsigned( 20,8)),
			9115 => std_logic_vector(to_unsigned( 199,8)),
			9116 => std_logic_vector(to_unsigned( 122,8)),
			9117 => std_logic_vector(to_unsigned( 161,8)),
			9118 => std_logic_vector(to_unsigned( 160,8)),
			9119 => std_logic_vector(to_unsigned( 191,8)),
			9120 => std_logic_vector(to_unsigned( 36,8)),
			9121 => std_logic_vector(to_unsigned( 183,8)),
			9122 => std_logic_vector(to_unsigned( 224,8)),
			9123 => std_logic_vector(to_unsigned( 49,8)),
			9124 => std_logic_vector(to_unsigned( 34,8)),
			9125 => std_logic_vector(to_unsigned( 113,8)),
			9126 => std_logic_vector(to_unsigned( 161,8)),
			9127 => std_logic_vector(to_unsigned( 116,8)),
			9128 => std_logic_vector(to_unsigned( 150,8)),
			9129 => std_logic_vector(to_unsigned( 2,8)),
			9130 => std_logic_vector(to_unsigned( 33,8)),
			9131 => std_logic_vector(to_unsigned( 172,8)),
			9132 => std_logic_vector(to_unsigned( 145,8)),
			9133 => std_logic_vector(to_unsigned( 56,8)),
			9134 => std_logic_vector(to_unsigned( 35,8)),
			9135 => std_logic_vector(to_unsigned( 111,8)),
			9136 => std_logic_vector(to_unsigned( 47,8)),
			9137 => std_logic_vector(to_unsigned( 46,8)),
			9138 => std_logic_vector(to_unsigned( 222,8)),
			9139 => std_logic_vector(to_unsigned( 170,8)),
			9140 => std_logic_vector(to_unsigned( 212,8)),
			9141 => std_logic_vector(to_unsigned( 53,8)),
			9142 => std_logic_vector(to_unsigned( 44,8)),
			9143 => std_logic_vector(to_unsigned( 130,8)),
			9144 => std_logic_vector(to_unsigned( 92,8)),
			9145 => std_logic_vector(to_unsigned( 134,8)),
			9146 => std_logic_vector(to_unsigned( 49,8)),
			9147 => std_logic_vector(to_unsigned( 169,8)),
			9148 => std_logic_vector(to_unsigned( 31,8)),
			9149 => std_logic_vector(to_unsigned( 131,8)),
			9150 => std_logic_vector(to_unsigned( 66,8)),
			9151 => std_logic_vector(to_unsigned( 122,8)),
			9152 => std_logic_vector(to_unsigned( 56,8)),
			9153 => std_logic_vector(to_unsigned( 222,8)),
			9154 => std_logic_vector(to_unsigned( 69,8)),
			9155 => std_logic_vector(to_unsigned( 147,8)),
			9156 => std_logic_vector(to_unsigned( 158,8)),
			9157 => std_logic_vector(to_unsigned( 248,8)),
			9158 => std_logic_vector(to_unsigned( 1,8)),
			9159 => std_logic_vector(to_unsigned( 49,8)),
			9160 => std_logic_vector(to_unsigned( 243,8)),
			9161 => std_logic_vector(to_unsigned( 16,8)),
			9162 => std_logic_vector(to_unsigned( 91,8)),
			9163 => std_logic_vector(to_unsigned( 36,8)),
			9164 => std_logic_vector(to_unsigned( 184,8)),
			9165 => std_logic_vector(to_unsigned( 24,8)),
			9166 => std_logic_vector(to_unsigned( 130,8)),
			9167 => std_logic_vector(to_unsigned( 46,8)),
			9168 => std_logic_vector(to_unsigned( 169,8)),
			9169 => std_logic_vector(to_unsigned( 79,8)),
			9170 => std_logic_vector(to_unsigned( 56,8)),
			9171 => std_logic_vector(to_unsigned( 102,8)),
			9172 => std_logic_vector(to_unsigned( 56,8)),
			9173 => std_logic_vector(to_unsigned( 161,8)),
			9174 => std_logic_vector(to_unsigned( 182,8)),
			9175 => std_logic_vector(to_unsigned( 132,8)),
			9176 => std_logic_vector(to_unsigned( 193,8)),
			9177 => std_logic_vector(to_unsigned( 119,8)),
			9178 => std_logic_vector(to_unsigned( 5,8)),
			9179 => std_logic_vector(to_unsigned( 159,8)),
			9180 => std_logic_vector(to_unsigned( 209,8)),
			9181 => std_logic_vector(to_unsigned( 233,8)),
			9182 => std_logic_vector(to_unsigned( 3,8)),
			9183 => std_logic_vector(to_unsigned( 150,8)),
			9184 => std_logic_vector(to_unsigned( 161,8)),
			9185 => std_logic_vector(to_unsigned( 82,8)),
			9186 => std_logic_vector(to_unsigned( 56,8)),
			9187 => std_logic_vector(to_unsigned( 139,8)),
			9188 => std_logic_vector(to_unsigned( 30,8)),
			9189 => std_logic_vector(to_unsigned( 123,8)),
			9190 => std_logic_vector(to_unsigned( 50,8)),
			9191 => std_logic_vector(to_unsigned( 88,8)),
			9192 => std_logic_vector(to_unsigned( 140,8)),
			9193 => std_logic_vector(to_unsigned( 80,8)),
			9194 => std_logic_vector(to_unsigned( 7,8)),
			9195 => std_logic_vector(to_unsigned( 210,8)),
			9196 => std_logic_vector(to_unsigned( 248,8)),
			9197 => std_logic_vector(to_unsigned( 51,8)),
			9198 => std_logic_vector(to_unsigned( 140,8)),
			9199 => std_logic_vector(to_unsigned( 29,8)),
			9200 => std_logic_vector(to_unsigned( 138,8)),
			9201 => std_logic_vector(to_unsigned( 247,8)),
			9202 => std_logic_vector(to_unsigned( 42,8)),
			9203 => std_logic_vector(to_unsigned( 157,8)),
			9204 => std_logic_vector(to_unsigned( 191,8)),
			9205 => std_logic_vector(to_unsigned( 65,8)),
			9206 => std_logic_vector(to_unsigned( 15,8)),
			9207 => std_logic_vector(to_unsigned( 109,8)),
			9208 => std_logic_vector(to_unsigned( 191,8)),
			9209 => std_logic_vector(to_unsigned( 153,8)),
			9210 => std_logic_vector(to_unsigned( 118,8)),
			9211 => std_logic_vector(to_unsigned( 160,8)),
			9212 => std_logic_vector(to_unsigned( 14,8)),
			9213 => std_logic_vector(to_unsigned( 123,8)),
			9214 => std_logic_vector(to_unsigned( 59,8)),
			9215 => std_logic_vector(to_unsigned( 185,8)),
			9216 => std_logic_vector(to_unsigned( 250,8)),
			9217 => std_logic_vector(to_unsigned( 250,8)),
			9218 => std_logic_vector(to_unsigned( 24,8)),
			9219 => std_logic_vector(to_unsigned( 71,8)),
			9220 => std_logic_vector(to_unsigned( 246,8)),
			9221 => std_logic_vector(to_unsigned( 190,8)),
			9222 => std_logic_vector(to_unsigned( 66,8)),
			9223 => std_logic_vector(to_unsigned( 186,8)),
			9224 => std_logic_vector(to_unsigned( 129,8)),
			9225 => std_logic_vector(to_unsigned( 229,8)),
			9226 => std_logic_vector(to_unsigned( 156,8)),
			9227 => std_logic_vector(to_unsigned( 39,8)),
			9228 => std_logic_vector(to_unsigned( 198,8)),
			9229 => std_logic_vector(to_unsigned( 91,8)),
			9230 => std_logic_vector(to_unsigned( 147,8)),
			9231 => std_logic_vector(to_unsigned( 160,8)),
			9232 => std_logic_vector(to_unsigned( 156,8)),
			9233 => std_logic_vector(to_unsigned( 222,8)),
			9234 => std_logic_vector(to_unsigned( 224,8)),
			9235 => std_logic_vector(to_unsigned( 232,8)),
			9236 => std_logic_vector(to_unsigned( 78,8)),
			9237 => std_logic_vector(to_unsigned( 188,8)),
			9238 => std_logic_vector(to_unsigned( 14,8)),
			9239 => std_logic_vector(to_unsigned( 4,8)),
			9240 => std_logic_vector(to_unsigned( 61,8)),
			9241 => std_logic_vector(to_unsigned( 11,8)),
			9242 => std_logic_vector(to_unsigned( 87,8)),
			9243 => std_logic_vector(to_unsigned( 92,8)),
			9244 => std_logic_vector(to_unsigned( 215,8)),
			9245 => std_logic_vector(to_unsigned( 3,8)),
			9246 => std_logic_vector(to_unsigned( 184,8)),
			9247 => std_logic_vector(to_unsigned( 93,8)),
			9248 => std_logic_vector(to_unsigned( 197,8)),
			9249 => std_logic_vector(to_unsigned( 93,8)),
			9250 => std_logic_vector(to_unsigned( 81,8)),
			9251 => std_logic_vector(to_unsigned( 205,8)),
			9252 => std_logic_vector(to_unsigned( 54,8)),
			9253 => std_logic_vector(to_unsigned( 185,8)),
			9254 => std_logic_vector(to_unsigned( 107,8)),
			9255 => std_logic_vector(to_unsigned( 38,8)),
			9256 => std_logic_vector(to_unsigned( 94,8)),
			9257 => std_logic_vector(to_unsigned( 80,8)),
			9258 => std_logic_vector(to_unsigned( 225,8)),
			9259 => std_logic_vector(to_unsigned( 55,8)),
			9260 => std_logic_vector(to_unsigned( 19,8)),
			9261 => std_logic_vector(to_unsigned( 121,8)),
			9262 => std_logic_vector(to_unsigned( 90,8)),
			9263 => std_logic_vector(to_unsigned( 29,8)),
			9264 => std_logic_vector(to_unsigned( 95,8)),
			9265 => std_logic_vector(to_unsigned( 172,8)),
			9266 => std_logic_vector(to_unsigned( 50,8)),
			9267 => std_logic_vector(to_unsigned( 7,8)),
			9268 => std_logic_vector(to_unsigned( 79,8)),
			9269 => std_logic_vector(to_unsigned( 101,8)),
			9270 => std_logic_vector(to_unsigned( 103,8)),
			9271 => std_logic_vector(to_unsigned( 18,8)),
			9272 => std_logic_vector(to_unsigned( 171,8)),
			9273 => std_logic_vector(to_unsigned( 90,8)),
			9274 => std_logic_vector(to_unsigned( 210,8)),
			9275 => std_logic_vector(to_unsigned( 1,8)),
			9276 => std_logic_vector(to_unsigned( 17,8)),
			9277 => std_logic_vector(to_unsigned( 147,8)),
			9278 => std_logic_vector(to_unsigned( 194,8)),
			9279 => std_logic_vector(to_unsigned( 228,8)),
			9280 => std_logic_vector(to_unsigned( 238,8)),
			9281 => std_logic_vector(to_unsigned( 232,8)),
			9282 => std_logic_vector(to_unsigned( 30,8)),
			9283 => std_logic_vector(to_unsigned( 16,8)),
			9284 => std_logic_vector(to_unsigned( 82,8)),
			9285 => std_logic_vector(to_unsigned( 122,8)),
			9286 => std_logic_vector(to_unsigned( 119,8)),
			9287 => std_logic_vector(to_unsigned( 149,8)),
			9288 => std_logic_vector(to_unsigned( 169,8)),
			9289 => std_logic_vector(to_unsigned( 91,8)),
			9290 => std_logic_vector(to_unsigned( 66,8)),
			9291 => std_logic_vector(to_unsigned( 44,8)),
			9292 => std_logic_vector(to_unsigned( 45,8)),
			9293 => std_logic_vector(to_unsigned( 248,8)),
			9294 => std_logic_vector(to_unsigned( 218,8)),
			9295 => std_logic_vector(to_unsigned( 25,8)),
			9296 => std_logic_vector(to_unsigned( 175,8)),
			9297 => std_logic_vector(to_unsigned( 224,8)),
			9298 => std_logic_vector(to_unsigned( 243,8)),
			9299 => std_logic_vector(to_unsigned( 23,8)),
			9300 => std_logic_vector(to_unsigned( 51,8)),
			9301 => std_logic_vector(to_unsigned( 131,8)),
			9302 => std_logic_vector(to_unsigned( 89,8)),
			9303 => std_logic_vector(to_unsigned( 239,8)),
			9304 => std_logic_vector(to_unsigned( 74,8)),
			9305 => std_logic_vector(to_unsigned( 146,8)),
			9306 => std_logic_vector(to_unsigned( 139,8)),
			9307 => std_logic_vector(to_unsigned( 123,8)),
			9308 => std_logic_vector(to_unsigned( 195,8)),
			9309 => std_logic_vector(to_unsigned( 2,8)),
			9310 => std_logic_vector(to_unsigned( 218,8)),
			9311 => std_logic_vector(to_unsigned( 56,8)),
			9312 => std_logic_vector(to_unsigned( 173,8)),
			9313 => std_logic_vector(to_unsigned( 127,8)),
			9314 => std_logic_vector(to_unsigned( 58,8)),
			9315 => std_logic_vector(to_unsigned( 6,8)),
			9316 => std_logic_vector(to_unsigned( 126,8)),
			9317 => std_logic_vector(to_unsigned( 22,8)),
			9318 => std_logic_vector(to_unsigned( 179,8)),
			9319 => std_logic_vector(to_unsigned( 111,8)),
			9320 => std_logic_vector(to_unsigned( 178,8)),
			9321 => std_logic_vector(to_unsigned( 104,8)),
			9322 => std_logic_vector(to_unsigned( 180,8)),
			9323 => std_logic_vector(to_unsigned( 70,8)),
			9324 => std_logic_vector(to_unsigned( 79,8)),
			9325 => std_logic_vector(to_unsigned( 125,8)),
			9326 => std_logic_vector(to_unsigned( 235,8)),
			9327 => std_logic_vector(to_unsigned( 244,8)),
			9328 => std_logic_vector(to_unsigned( 248,8)),
			9329 => std_logic_vector(to_unsigned( 233,8)),
			9330 => std_logic_vector(to_unsigned( 209,8)),
			9331 => std_logic_vector(to_unsigned( 32,8)),
			9332 => std_logic_vector(to_unsigned( 207,8)),
			9333 => std_logic_vector(to_unsigned( 216,8)),
			9334 => std_logic_vector(to_unsigned( 151,8)),
			9335 => std_logic_vector(to_unsigned( 160,8)),
			9336 => std_logic_vector(to_unsigned( 35,8)),
			9337 => std_logic_vector(to_unsigned( 84,8)),
			9338 => std_logic_vector(to_unsigned( 80,8)),
			9339 => std_logic_vector(to_unsigned( 142,8)),
			9340 => std_logic_vector(to_unsigned( 37,8)),
			9341 => std_logic_vector(to_unsigned( 240,8)),
			9342 => std_logic_vector(to_unsigned( 123,8)),
			9343 => std_logic_vector(to_unsigned( 156,8)),
			9344 => std_logic_vector(to_unsigned( 144,8)),
			9345 => std_logic_vector(to_unsigned( 204,8)),
			9346 => std_logic_vector(to_unsigned( 99,8)),
			9347 => std_logic_vector(to_unsigned( 217,8)),
			9348 => std_logic_vector(to_unsigned( 74,8)),
			9349 => std_logic_vector(to_unsigned( 88,8)),
			9350 => std_logic_vector(to_unsigned( 176,8)),
			9351 => std_logic_vector(to_unsigned( 46,8)),
			9352 => std_logic_vector(to_unsigned( 52,8)),
			9353 => std_logic_vector(to_unsigned( 23,8)),
			9354 => std_logic_vector(to_unsigned( 81,8)),
			9355 => std_logic_vector(to_unsigned( 175,8)),
			9356 => std_logic_vector(to_unsigned( 123,8)),
			9357 => std_logic_vector(to_unsigned( 206,8)),
			9358 => std_logic_vector(to_unsigned( 77,8)),
			9359 => std_logic_vector(to_unsigned( 121,8)),
			9360 => std_logic_vector(to_unsigned( 222,8)),
			9361 => std_logic_vector(to_unsigned( 97,8)),
			9362 => std_logic_vector(to_unsigned( 236,8)),
			9363 => std_logic_vector(to_unsigned( 66,8)),
			9364 => std_logic_vector(to_unsigned( 254,8)),
			9365 => std_logic_vector(to_unsigned( 127,8)),
			9366 => std_logic_vector(to_unsigned( 12,8)),
			9367 => std_logic_vector(to_unsigned( 43,8)),
			9368 => std_logic_vector(to_unsigned( 206,8)),
			9369 => std_logic_vector(to_unsigned( 31,8)),
			9370 => std_logic_vector(to_unsigned( 141,8)),
			9371 => std_logic_vector(to_unsigned( 145,8)),
			9372 => std_logic_vector(to_unsigned( 107,8)),
			9373 => std_logic_vector(to_unsigned( 188,8)),
			9374 => std_logic_vector(to_unsigned( 163,8)),
			9375 => std_logic_vector(to_unsigned( 247,8)),
			9376 => std_logic_vector(to_unsigned( 162,8)),
			9377 => std_logic_vector(to_unsigned( 222,8)),
			9378 => std_logic_vector(to_unsigned( 228,8)),
			9379 => std_logic_vector(to_unsigned( 41,8)),
			9380 => std_logic_vector(to_unsigned( 127,8)),
			9381 => std_logic_vector(to_unsigned( 231,8)),
			9382 => std_logic_vector(to_unsigned( 90,8)),
			9383 => std_logic_vector(to_unsigned( 96,8)),
			9384 => std_logic_vector(to_unsigned( 8,8)),
			9385 => std_logic_vector(to_unsigned( 72,8)),
			9386 => std_logic_vector(to_unsigned( 129,8)),
			9387 => std_logic_vector(to_unsigned( 7,8)),
			9388 => std_logic_vector(to_unsigned( 33,8)),
			9389 => std_logic_vector(to_unsigned( 117,8)),
			9390 => std_logic_vector(to_unsigned( 52,8)),
			9391 => std_logic_vector(to_unsigned( 0,8)),
			9392 => std_logic_vector(to_unsigned( 202,8)),
			9393 => std_logic_vector(to_unsigned( 196,8)),
			9394 => std_logic_vector(to_unsigned( 193,8)),
			9395 => std_logic_vector(to_unsigned( 147,8)),
			9396 => std_logic_vector(to_unsigned( 209,8)),
			9397 => std_logic_vector(to_unsigned( 16,8)),
			9398 => std_logic_vector(to_unsigned( 140,8)),
			9399 => std_logic_vector(to_unsigned( 108,8)),
			9400 => std_logic_vector(to_unsigned( 18,8)),
			9401 => std_logic_vector(to_unsigned( 235,8)),
			9402 => std_logic_vector(to_unsigned( 210,8)),
			9403 => std_logic_vector(to_unsigned( 56,8)),
			9404 => std_logic_vector(to_unsigned( 5,8)),
			9405 => std_logic_vector(to_unsigned( 110,8)),
			9406 => std_logic_vector(to_unsigned( 121,8)),
			9407 => std_logic_vector(to_unsigned( 156,8)),
			9408 => std_logic_vector(to_unsigned( 127,8)),
			9409 => std_logic_vector(to_unsigned( 236,8)),
			9410 => std_logic_vector(to_unsigned( 115,8)),
			9411 => std_logic_vector(to_unsigned( 83,8)),
			9412 => std_logic_vector(to_unsigned( 6,8)),
			9413 => std_logic_vector(to_unsigned( 228,8)),
			9414 => std_logic_vector(to_unsigned( 82,8)),
			9415 => std_logic_vector(to_unsigned( 168,8)),
			9416 => std_logic_vector(to_unsigned( 35,8)),
			9417 => std_logic_vector(to_unsigned( 17,8)),
			9418 => std_logic_vector(to_unsigned( 7,8)),
			9419 => std_logic_vector(to_unsigned( 138,8)),
			9420 => std_logic_vector(to_unsigned( 166,8)),
			9421 => std_logic_vector(to_unsigned( 95,8)),
			9422 => std_logic_vector(to_unsigned( 5,8)),
			9423 => std_logic_vector(to_unsigned( 87,8)),
			9424 => std_logic_vector(to_unsigned( 18,8)),
			9425 => std_logic_vector(to_unsigned( 115,8)),
			9426 => std_logic_vector(to_unsigned( 150,8)),
			9427 => std_logic_vector(to_unsigned( 96,8)),
			9428 => std_logic_vector(to_unsigned( 145,8)),
			9429 => std_logic_vector(to_unsigned( 239,8)),
			9430 => std_logic_vector(to_unsigned( 104,8)),
			9431 => std_logic_vector(to_unsigned( 52,8)),
			9432 => std_logic_vector(to_unsigned( 6,8)),
			9433 => std_logic_vector(to_unsigned( 166,8)),
			9434 => std_logic_vector(to_unsigned( 55,8)),
			9435 => std_logic_vector(to_unsigned( 188,8)),
			9436 => std_logic_vector(to_unsigned( 118,8)),
			9437 => std_logic_vector(to_unsigned( 177,8)),
			9438 => std_logic_vector(to_unsigned( 6,8)),
			9439 => std_logic_vector(to_unsigned( 243,8)),
			9440 => std_logic_vector(to_unsigned( 246,8)),
			9441 => std_logic_vector(to_unsigned( 10,8)),
			9442 => std_logic_vector(to_unsigned( 14,8)),
			9443 => std_logic_vector(to_unsigned( 17,8)),
			9444 => std_logic_vector(to_unsigned( 168,8)),
			9445 => std_logic_vector(to_unsigned( 34,8)),
			9446 => std_logic_vector(to_unsigned( 140,8)),
			9447 => std_logic_vector(to_unsigned( 132,8)),
			9448 => std_logic_vector(to_unsigned( 143,8)),
			9449 => std_logic_vector(to_unsigned( 122,8)),
			9450 => std_logic_vector(to_unsigned( 75,8)),
			9451 => std_logic_vector(to_unsigned( 217,8)),
			9452 => std_logic_vector(to_unsigned( 225,8)),
			9453 => std_logic_vector(to_unsigned( 227,8)),
			9454 => std_logic_vector(to_unsigned( 214,8)),
			9455 => std_logic_vector(to_unsigned( 10,8)),
			9456 => std_logic_vector(to_unsigned( 151,8)),
			9457 => std_logic_vector(to_unsigned( 245,8)),
			9458 => std_logic_vector(to_unsigned( 216,8)),
			9459 => std_logic_vector(to_unsigned( 108,8)),
			9460 => std_logic_vector(to_unsigned( 114,8)),
			9461 => std_logic_vector(to_unsigned( 45,8)),
			9462 => std_logic_vector(to_unsigned( 245,8)),
			9463 => std_logic_vector(to_unsigned( 59,8)),
			9464 => std_logic_vector(to_unsigned( 1,8)),
			9465 => std_logic_vector(to_unsigned( 165,8)),
			9466 => std_logic_vector(to_unsigned( 23,8)),
			9467 => std_logic_vector(to_unsigned( 23,8)),
			9468 => std_logic_vector(to_unsigned( 55,8)),
			9469 => std_logic_vector(to_unsigned( 221,8)),
			9470 => std_logic_vector(to_unsigned( 86,8)),
			9471 => std_logic_vector(to_unsigned( 102,8)),
			9472 => std_logic_vector(to_unsigned( 60,8)),
			9473 => std_logic_vector(to_unsigned( 109,8)),
			9474 => std_logic_vector(to_unsigned( 125,8)),
			9475 => std_logic_vector(to_unsigned( 100,8)),
			9476 => std_logic_vector(to_unsigned( 108,8)),
			9477 => std_logic_vector(to_unsigned( 101,8)),
			9478 => std_logic_vector(to_unsigned( 250,8)),
			9479 => std_logic_vector(to_unsigned( 71,8)),
			9480 => std_logic_vector(to_unsigned( 154,8)),
			9481 => std_logic_vector(to_unsigned( 55,8)),
			9482 => std_logic_vector(to_unsigned( 93,8)),
			9483 => std_logic_vector(to_unsigned( 82,8)),
			9484 => std_logic_vector(to_unsigned( 212,8)),
			9485 => std_logic_vector(to_unsigned( 123,8)),
			9486 => std_logic_vector(to_unsigned( 207,8)),
			9487 => std_logic_vector(to_unsigned( 140,8)),
			9488 => std_logic_vector(to_unsigned( 73,8)),
			9489 => std_logic_vector(to_unsigned( 174,8)),
			9490 => std_logic_vector(to_unsigned( 146,8)),
			9491 => std_logic_vector(to_unsigned( 215,8)),
			9492 => std_logic_vector(to_unsigned( 97,8)),
			9493 => std_logic_vector(to_unsigned( 96,8)),
			9494 => std_logic_vector(to_unsigned( 196,8)),
			9495 => std_logic_vector(to_unsigned( 103,8)),
			9496 => std_logic_vector(to_unsigned( 136,8)),
			9497 => std_logic_vector(to_unsigned( 85,8)),
			9498 => std_logic_vector(to_unsigned( 212,8)),
			9499 => std_logic_vector(to_unsigned( 23,8)),
			9500 => std_logic_vector(to_unsigned( 77,8)),
			9501 => std_logic_vector(to_unsigned( 239,8)),
			9502 => std_logic_vector(to_unsigned( 18,8)),
			9503 => std_logic_vector(to_unsigned( 162,8)),
			9504 => std_logic_vector(to_unsigned( 249,8)),
			9505 => std_logic_vector(to_unsigned( 53,8)),
			9506 => std_logic_vector(to_unsigned( 212,8)),
			9507 => std_logic_vector(to_unsigned( 246,8)),
			9508 => std_logic_vector(to_unsigned( 81,8)),
			9509 => std_logic_vector(to_unsigned( 211,8)),
			9510 => std_logic_vector(to_unsigned( 91,8)),
			9511 => std_logic_vector(to_unsigned( 177,8)),
			9512 => std_logic_vector(to_unsigned( 248,8)),
			9513 => std_logic_vector(to_unsigned( 70,8)),
			9514 => std_logic_vector(to_unsigned( 173,8)),
			9515 => std_logic_vector(to_unsigned( 108,8)),
			9516 => std_logic_vector(to_unsigned( 195,8)),
			9517 => std_logic_vector(to_unsigned( 46,8)),
			9518 => std_logic_vector(to_unsigned( 119,8)),
			9519 => std_logic_vector(to_unsigned( 16,8)),
			9520 => std_logic_vector(to_unsigned( 152,8)),
			9521 => std_logic_vector(to_unsigned( 53,8)),
			9522 => std_logic_vector(to_unsigned( 223,8)),
			9523 => std_logic_vector(to_unsigned( 233,8)),
			9524 => std_logic_vector(to_unsigned( 190,8)),
			9525 => std_logic_vector(to_unsigned( 232,8)),
			9526 => std_logic_vector(to_unsigned( 198,8)),
			9527 => std_logic_vector(to_unsigned( 161,8)),
			9528 => std_logic_vector(to_unsigned( 219,8)),
			9529 => std_logic_vector(to_unsigned( 24,8)),
			9530 => std_logic_vector(to_unsigned( 169,8)),
			9531 => std_logic_vector(to_unsigned( 16,8)),
			9532 => std_logic_vector(to_unsigned( 139,8)),
			9533 => std_logic_vector(to_unsigned( 35,8)),
			9534 => std_logic_vector(to_unsigned( 141,8)),
			9535 => std_logic_vector(to_unsigned( 145,8)),
			9536 => std_logic_vector(to_unsigned( 157,8)),
			9537 => std_logic_vector(to_unsigned( 26,8)),
			9538 => std_logic_vector(to_unsigned( 221,8)),
			9539 => std_logic_vector(to_unsigned( 73,8)),
			9540 => std_logic_vector(to_unsigned( 0,8)),
			9541 => std_logic_vector(to_unsigned( 162,8)),
			9542 => std_logic_vector(to_unsigned( 23,8)),
			9543 => std_logic_vector(to_unsigned( 238,8)),
			9544 => std_logic_vector(to_unsigned( 127,8)),
			9545 => std_logic_vector(to_unsigned( 77,8)),
			9546 => std_logic_vector(to_unsigned( 40,8)),
			9547 => std_logic_vector(to_unsigned( 54,8)),
			9548 => std_logic_vector(to_unsigned( 53,8)),
			9549 => std_logic_vector(to_unsigned( 160,8)),
			9550 => std_logic_vector(to_unsigned( 226,8)),
			9551 => std_logic_vector(to_unsigned( 240,8)),
			9552 => std_logic_vector(to_unsigned( 173,8)),
			9553 => std_logic_vector(to_unsigned( 116,8)),
			9554 => std_logic_vector(to_unsigned( 56,8)),
			9555 => std_logic_vector(to_unsigned( 234,8)),
			9556 => std_logic_vector(to_unsigned( 46,8)),
			9557 => std_logic_vector(to_unsigned( 180,8)),
			9558 => std_logic_vector(to_unsigned( 248,8)),
			9559 => std_logic_vector(to_unsigned( 187,8)),
			9560 => std_logic_vector(to_unsigned( 249,8)),
			9561 => std_logic_vector(to_unsigned( 102,8)),
			9562 => std_logic_vector(to_unsigned( 252,8)),
			9563 => std_logic_vector(to_unsigned( 27,8)),
			9564 => std_logic_vector(to_unsigned( 36,8)),
			9565 => std_logic_vector(to_unsigned( 169,8)),
			9566 => std_logic_vector(to_unsigned( 209,8)),
			9567 => std_logic_vector(to_unsigned( 151,8)),
			9568 => std_logic_vector(to_unsigned( 231,8)),
			9569 => std_logic_vector(to_unsigned( 29,8)),
			9570 => std_logic_vector(to_unsigned( 235,8)),
			9571 => std_logic_vector(to_unsigned( 135,8)),
			9572 => std_logic_vector(to_unsigned( 151,8)),
			9573 => std_logic_vector(to_unsigned( 147,8)),
			9574 => std_logic_vector(to_unsigned( 25,8)),
			9575 => std_logic_vector(to_unsigned( 79,8)),
			9576 => std_logic_vector(to_unsigned( 193,8)),
			9577 => std_logic_vector(to_unsigned( 70,8)),
			9578 => std_logic_vector(to_unsigned( 62,8)),
			9579 => std_logic_vector(to_unsigned( 246,8)),
			9580 => std_logic_vector(to_unsigned( 64,8)),
			9581 => std_logic_vector(to_unsigned( 43,8)),
			9582 => std_logic_vector(to_unsigned( 158,8)),
			9583 => std_logic_vector(to_unsigned( 175,8)),
			9584 => std_logic_vector(to_unsigned( 71,8)),
			9585 => std_logic_vector(to_unsigned( 232,8)),
			9586 => std_logic_vector(to_unsigned( 239,8)),
			9587 => std_logic_vector(to_unsigned( 44,8)),
			9588 => std_logic_vector(to_unsigned( 177,8)),
			9589 => std_logic_vector(to_unsigned( 212,8)),
			9590 => std_logic_vector(to_unsigned( 72,8)),
			9591 => std_logic_vector(to_unsigned( 131,8)),
			9592 => std_logic_vector(to_unsigned( 13,8)),
			9593 => std_logic_vector(to_unsigned( 11,8)),
			9594 => std_logic_vector(to_unsigned( 71,8)),
			9595 => std_logic_vector(to_unsigned( 41,8)),
			9596 => std_logic_vector(to_unsigned( 130,8)),
			9597 => std_logic_vector(to_unsigned( 197,8)),
			9598 => std_logic_vector(to_unsigned( 205,8)),
			9599 => std_logic_vector(to_unsigned( 166,8)),
			9600 => std_logic_vector(to_unsigned( 216,8)),
			9601 => std_logic_vector(to_unsigned( 183,8)),
			9602 => std_logic_vector(to_unsigned( 38,8)),
			9603 => std_logic_vector(to_unsigned( 85,8)),
			9604 => std_logic_vector(to_unsigned( 146,8)),
			9605 => std_logic_vector(to_unsigned( 53,8)),
			9606 => std_logic_vector(to_unsigned( 124,8)),
			9607 => std_logic_vector(to_unsigned( 118,8)),
			9608 => std_logic_vector(to_unsigned( 188,8)),
			9609 => std_logic_vector(to_unsigned( 151,8)),
			9610 => std_logic_vector(to_unsigned( 103,8)),
			9611 => std_logic_vector(to_unsigned( 101,8)),
			9612 => std_logic_vector(to_unsigned( 106,8)),
			9613 => std_logic_vector(to_unsigned( 48,8)),
			9614 => std_logic_vector(to_unsigned( 60,8)),
			9615 => std_logic_vector(to_unsigned( 199,8)),
			9616 => std_logic_vector(to_unsigned( 170,8)),
			9617 => std_logic_vector(to_unsigned( 167,8)),
			9618 => std_logic_vector(to_unsigned( 159,8)),
			9619 => std_logic_vector(to_unsigned( 188,8)),
			9620 => std_logic_vector(to_unsigned( 228,8)),
			9621 => std_logic_vector(to_unsigned( 183,8)),
			9622 => std_logic_vector(to_unsigned( 211,8)),
			9623 => std_logic_vector(to_unsigned( 250,8)),
			9624 => std_logic_vector(to_unsigned( 34,8)),
			9625 => std_logic_vector(to_unsigned( 228,8)),
			9626 => std_logic_vector(to_unsigned( 8,8)),
			9627 => std_logic_vector(to_unsigned( 28,8)),
			9628 => std_logic_vector(to_unsigned( 99,8)),
			9629 => std_logic_vector(to_unsigned( 122,8)),
			9630 => std_logic_vector(to_unsigned( 146,8)),
			9631 => std_logic_vector(to_unsigned( 172,8)),
			9632 => std_logic_vector(to_unsigned( 212,8)),
			9633 => std_logic_vector(to_unsigned( 87,8)),
			9634 => std_logic_vector(to_unsigned( 231,8)),
			9635 => std_logic_vector(to_unsigned( 43,8)),
			9636 => std_logic_vector(to_unsigned( 145,8)),
			9637 => std_logic_vector(to_unsigned( 241,8)),
			9638 => std_logic_vector(to_unsigned( 166,8)),
			9639 => std_logic_vector(to_unsigned( 48,8)),
			9640 => std_logic_vector(to_unsigned( 34,8)),
			9641 => std_logic_vector(to_unsigned( 44,8)),
			9642 => std_logic_vector(to_unsigned( 40,8)),
			9643 => std_logic_vector(to_unsigned( 234,8)),
			9644 => std_logic_vector(to_unsigned( 201,8)),
			9645 => std_logic_vector(to_unsigned( 164,8)),
			9646 => std_logic_vector(to_unsigned( 134,8)),
			9647 => std_logic_vector(to_unsigned( 172,8)),
			9648 => std_logic_vector(to_unsigned( 142,8)),
			9649 => std_logic_vector(to_unsigned( 119,8)),
			9650 => std_logic_vector(to_unsigned( 162,8)),
			9651 => std_logic_vector(to_unsigned( 43,8)),
			9652 => std_logic_vector(to_unsigned( 241,8)),
			9653 => std_logic_vector(to_unsigned( 99,8)),
			9654 => std_logic_vector(to_unsigned( 142,8)),
			9655 => std_logic_vector(to_unsigned( 173,8)),
			9656 => std_logic_vector(to_unsigned( 222,8)),
			9657 => std_logic_vector(to_unsigned( 128,8)),
			9658 => std_logic_vector(to_unsigned( 196,8)),
			9659 => std_logic_vector(to_unsigned( 225,8)),
			9660 => std_logic_vector(to_unsigned( 223,8)),
			9661 => std_logic_vector(to_unsigned( 114,8)),
			9662 => std_logic_vector(to_unsigned( 208,8)),
			9663 => std_logic_vector(to_unsigned( 134,8)),
			9664 => std_logic_vector(to_unsigned( 155,8)),
			9665 => std_logic_vector(to_unsigned( 42,8)),
			9666 => std_logic_vector(to_unsigned( 3,8)),
			9667 => std_logic_vector(to_unsigned( 205,8)),
			9668 => std_logic_vector(to_unsigned( 49,8)),
			9669 => std_logic_vector(to_unsigned( 13,8)),
			9670 => std_logic_vector(to_unsigned( 250,8)),
			9671 => std_logic_vector(to_unsigned( 150,8)),
			9672 => std_logic_vector(to_unsigned( 78,8)),
			9673 => std_logic_vector(to_unsigned( 163,8)),
			9674 => std_logic_vector(to_unsigned( 103,8)),
			9675 => std_logic_vector(to_unsigned( 137,8)),
			9676 => std_logic_vector(to_unsigned( 4,8)),
			9677 => std_logic_vector(to_unsigned( 156,8)),
			9678 => std_logic_vector(to_unsigned( 167,8)),
			9679 => std_logic_vector(to_unsigned( 145,8)),
			9680 => std_logic_vector(to_unsigned( 77,8)),
			9681 => std_logic_vector(to_unsigned( 163,8)),
			9682 => std_logic_vector(to_unsigned( 103,8)),
			9683 => std_logic_vector(to_unsigned( 252,8)),
			9684 => std_logic_vector(to_unsigned( 163,8)),
			9685 => std_logic_vector(to_unsigned( 58,8)),
			9686 => std_logic_vector(to_unsigned( 196,8)),
			9687 => std_logic_vector(to_unsigned( 231,8)),
			9688 => std_logic_vector(to_unsigned( 89,8)),
			9689 => std_logic_vector(to_unsigned( 59,8)),
			9690 => std_logic_vector(to_unsigned( 210,8)),
			9691 => std_logic_vector(to_unsigned( 232,8)),
			9692 => std_logic_vector(to_unsigned( 242,8)),
			9693 => std_logic_vector(to_unsigned( 37,8)),
			9694 => std_logic_vector(to_unsigned( 35,8)),
			9695 => std_logic_vector(to_unsigned( 215,8)),
			9696 => std_logic_vector(to_unsigned( 203,8)),
			9697 => std_logic_vector(to_unsigned( 89,8)),
			9698 => std_logic_vector(to_unsigned( 100,8)),
			9699 => std_logic_vector(to_unsigned( 183,8)),
			9700 => std_logic_vector(to_unsigned( 19,8)),
			9701 => std_logic_vector(to_unsigned( 164,8)),
			9702 => std_logic_vector(to_unsigned( 1,8)),
			9703 => std_logic_vector(to_unsigned( 23,8)),
			9704 => std_logic_vector(to_unsigned( 22,8)),
			9705 => std_logic_vector(to_unsigned( 94,8)),
			9706 => std_logic_vector(to_unsigned( 203,8)),
			9707 => std_logic_vector(to_unsigned( 121,8)),
			9708 => std_logic_vector(to_unsigned( 138,8)),
			9709 => std_logic_vector(to_unsigned( 127,8)),
			9710 => std_logic_vector(to_unsigned( 50,8)),
			9711 => std_logic_vector(to_unsigned( 77,8)),
			9712 => std_logic_vector(to_unsigned( 31,8)),
			9713 => std_logic_vector(to_unsigned( 83,8)),
			9714 => std_logic_vector(to_unsigned( 173,8)),
			9715 => std_logic_vector(to_unsigned( 84,8)),
			9716 => std_logic_vector(to_unsigned( 69,8)),
			9717 => std_logic_vector(to_unsigned( 211,8)),
			9718 => std_logic_vector(to_unsigned( 213,8)),
			9719 => std_logic_vector(to_unsigned( 32,8)),
			9720 => std_logic_vector(to_unsigned( 45,8)),
			9721 => std_logic_vector(to_unsigned( 115,8)),
			9722 => std_logic_vector(to_unsigned( 235,8)),
			9723 => std_logic_vector(to_unsigned( 96,8)),
			9724 => std_logic_vector(to_unsigned( 36,8)),
			9725 => std_logic_vector(to_unsigned( 11,8)),
			9726 => std_logic_vector(to_unsigned( 38,8)),
			9727 => std_logic_vector(to_unsigned( 92,8)),
			9728 => std_logic_vector(to_unsigned( 122,8)),
			9729 => std_logic_vector(to_unsigned( 197,8)),
			9730 => std_logic_vector(to_unsigned( 82,8)),
			9731 => std_logic_vector(to_unsigned( 21,8)),
			9732 => std_logic_vector(to_unsigned( 23,8)),
			9733 => std_logic_vector(to_unsigned( 178,8)),
			9734 => std_logic_vector(to_unsigned( 38,8)),
			9735 => std_logic_vector(to_unsigned( 216,8)),
			9736 => std_logic_vector(to_unsigned( 134,8)),
			9737 => std_logic_vector(to_unsigned( 123,8)),
			9738 => std_logic_vector(to_unsigned( 87,8)),
			9739 => std_logic_vector(to_unsigned( 9,8)),
			9740 => std_logic_vector(to_unsigned( 124,8)),
			9741 => std_logic_vector(to_unsigned( 121,8)),
			9742 => std_logic_vector(to_unsigned( 41,8)),
			9743 => std_logic_vector(to_unsigned( 40,8)),
			9744 => std_logic_vector(to_unsigned( 195,8)),
			9745 => std_logic_vector(to_unsigned( 189,8)),
			9746 => std_logic_vector(to_unsigned( 202,8)),
			9747 => std_logic_vector(to_unsigned( 130,8)),
			9748 => std_logic_vector(to_unsigned( 82,8)),
			9749 => std_logic_vector(to_unsigned( 160,8)),
			9750 => std_logic_vector(to_unsigned( 107,8)),
			9751 => std_logic_vector(to_unsigned( 21,8)),
			9752 => std_logic_vector(to_unsigned( 159,8)),
			9753 => std_logic_vector(to_unsigned( 4,8)),
			9754 => std_logic_vector(to_unsigned( 136,8)),
			9755 => std_logic_vector(to_unsigned( 222,8)),
			9756 => std_logic_vector(to_unsigned( 180,8)),
			9757 => std_logic_vector(to_unsigned( 107,8)),
			9758 => std_logic_vector(to_unsigned( 99,8)),
			9759 => std_logic_vector(to_unsigned( 104,8)),
			9760 => std_logic_vector(to_unsigned( 146,8)),
			9761 => std_logic_vector(to_unsigned( 253,8)),
			9762 => std_logic_vector(to_unsigned( 184,8)),
			9763 => std_logic_vector(to_unsigned( 60,8)),
			9764 => std_logic_vector(to_unsigned( 35,8)),
			9765 => std_logic_vector(to_unsigned( 0,8)),
			9766 => std_logic_vector(to_unsigned( 233,8)),
			9767 => std_logic_vector(to_unsigned( 108,8)),
			9768 => std_logic_vector(to_unsigned( 232,8)),
			9769 => std_logic_vector(to_unsigned( 196,8)),
			9770 => std_logic_vector(to_unsigned( 63,8)),
			9771 => std_logic_vector(to_unsigned( 56,8)),
			9772 => std_logic_vector(to_unsigned( 59,8)),
			9773 => std_logic_vector(to_unsigned( 20,8)),
			9774 => std_logic_vector(to_unsigned( 57,8)),
			9775 => std_logic_vector(to_unsigned( 237,8)),
			9776 => std_logic_vector(to_unsigned( 174,8)),
			9777 => std_logic_vector(to_unsigned( 137,8)),
			9778 => std_logic_vector(to_unsigned( 0,8)),
			9779 => std_logic_vector(to_unsigned( 48,8)),
			9780 => std_logic_vector(to_unsigned( 129,8)),
			9781 => std_logic_vector(to_unsigned( 75,8)),
			9782 => std_logic_vector(to_unsigned( 241,8)),
			9783 => std_logic_vector(to_unsigned( 151,8)),
			9784 => std_logic_vector(to_unsigned( 252,8)),
			9785 => std_logic_vector(to_unsigned( 27,8)),
			9786 => std_logic_vector(to_unsigned( 136,8)),
			9787 => std_logic_vector(to_unsigned( 220,8)),
			9788 => std_logic_vector(to_unsigned( 149,8)),
			9789 => std_logic_vector(to_unsigned( 16,8)),
			9790 => std_logic_vector(to_unsigned( 153,8)),
			9791 => std_logic_vector(to_unsigned( 11,8)),
			9792 => std_logic_vector(to_unsigned( 76,8)),
			9793 => std_logic_vector(to_unsigned( 229,8)),
			9794 => std_logic_vector(to_unsigned( 166,8)),
			9795 => std_logic_vector(to_unsigned( 141,8)),
			9796 => std_logic_vector(to_unsigned( 245,8)),
			9797 => std_logic_vector(to_unsigned( 134,8)),
			9798 => std_logic_vector(to_unsigned( 135,8)),
			9799 => std_logic_vector(to_unsigned( 8,8)),
			9800 => std_logic_vector(to_unsigned( 227,8)),
			9801 => std_logic_vector(to_unsigned( 137,8)),
			9802 => std_logic_vector(to_unsigned( 25,8)),
			9803 => std_logic_vector(to_unsigned( 27,8)),
			9804 => std_logic_vector(to_unsigned( 164,8)),
			9805 => std_logic_vector(to_unsigned( 198,8)),
			9806 => std_logic_vector(to_unsigned( 22,8)),
			9807 => std_logic_vector(to_unsigned( 41,8)),
			9808 => std_logic_vector(to_unsigned( 70,8)),
			9809 => std_logic_vector(to_unsigned( 194,8)),
			9810 => std_logic_vector(to_unsigned( 197,8)),
			9811 => std_logic_vector(to_unsigned( 127,8)),
			9812 => std_logic_vector(to_unsigned( 191,8)),
			9813 => std_logic_vector(to_unsigned( 23,8)),
			9814 => std_logic_vector(to_unsigned( 56,8)),
			9815 => std_logic_vector(to_unsigned( 245,8)),
			9816 => std_logic_vector(to_unsigned( 200,8)),
			9817 => std_logic_vector(to_unsigned( 33,8)),
			9818 => std_logic_vector(to_unsigned( 25,8)),
			9819 => std_logic_vector(to_unsigned( 100,8)),
			9820 => std_logic_vector(to_unsigned( 23,8)),
			9821 => std_logic_vector(to_unsigned( 153,8)),
			9822 => std_logic_vector(to_unsigned( 253,8)),
			9823 => std_logic_vector(to_unsigned( 29,8)),
			9824 => std_logic_vector(to_unsigned( 82,8)),
			9825 => std_logic_vector(to_unsigned( 76,8)),
			9826 => std_logic_vector(to_unsigned( 87,8)),
			9827 => std_logic_vector(to_unsigned( 1,8)),
			9828 => std_logic_vector(to_unsigned( 5,8)),
			9829 => std_logic_vector(to_unsigned( 50,8)),
			9830 => std_logic_vector(to_unsigned( 13,8)),
			9831 => std_logic_vector(to_unsigned( 75,8)),
			9832 => std_logic_vector(to_unsigned( 150,8)),
			9833 => std_logic_vector(to_unsigned( 67,8)),
			9834 => std_logic_vector(to_unsigned( 104,8)),
			9835 => std_logic_vector(to_unsigned( 13,8)),
			9836 => std_logic_vector(to_unsigned( 211,8)),
			9837 => std_logic_vector(to_unsigned( 15,8)),
			9838 => std_logic_vector(to_unsigned( 66,8)),
			9839 => std_logic_vector(to_unsigned( 224,8)),
			9840 => std_logic_vector(to_unsigned( 187,8)),
			9841 => std_logic_vector(to_unsigned( 211,8)),
			9842 => std_logic_vector(to_unsigned( 60,8)),
			9843 => std_logic_vector(to_unsigned( 178,8)),
			9844 => std_logic_vector(to_unsigned( 232,8)),
			9845 => std_logic_vector(to_unsigned( 197,8)),
			9846 => std_logic_vector(to_unsigned( 196,8)),
			9847 => std_logic_vector(to_unsigned( 219,8)),
			9848 => std_logic_vector(to_unsigned( 66,8)),
			9849 => std_logic_vector(to_unsigned( 52,8)),
			9850 => std_logic_vector(to_unsigned( 114,8)),
			9851 => std_logic_vector(to_unsigned( 60,8)),
			9852 => std_logic_vector(to_unsigned( 115,8)),
			9853 => std_logic_vector(to_unsigned( 191,8)),
			9854 => std_logic_vector(to_unsigned( 61,8)),
			9855 => std_logic_vector(to_unsigned( 216,8)),
			9856 => std_logic_vector(to_unsigned( 3,8)),
			9857 => std_logic_vector(to_unsigned( 129,8)),
			9858 => std_logic_vector(to_unsigned( 152,8)),
			9859 => std_logic_vector(to_unsigned( 131,8)),
			9860 => std_logic_vector(to_unsigned( 115,8)),
			9861 => std_logic_vector(to_unsigned( 254,8)),
			9862 => std_logic_vector(to_unsigned( 84,8)),
			9863 => std_logic_vector(to_unsigned( 151,8)),
			9864 => std_logic_vector(to_unsigned( 118,8)),
			9865 => std_logic_vector(to_unsigned( 79,8)),
			9866 => std_logic_vector(to_unsigned( 146,8)),
			9867 => std_logic_vector(to_unsigned( 239,8)),
			9868 => std_logic_vector(to_unsigned( 181,8)),
			9869 => std_logic_vector(to_unsigned( 188,8)),
			9870 => std_logic_vector(to_unsigned( 38,8)),
			9871 => std_logic_vector(to_unsigned( 119,8)),
			9872 => std_logic_vector(to_unsigned( 193,8)),
			9873 => std_logic_vector(to_unsigned( 45,8)),
			9874 => std_logic_vector(to_unsigned( 37,8)),
			9875 => std_logic_vector(to_unsigned( 34,8)),
			9876 => std_logic_vector(to_unsigned( 73,8)),
			9877 => std_logic_vector(to_unsigned( 197,8)),
			9878 => std_logic_vector(to_unsigned( 116,8)),
			9879 => std_logic_vector(to_unsigned( 109,8)),
			9880 => std_logic_vector(to_unsigned( 97,8)),
			9881 => std_logic_vector(to_unsigned( 163,8)),
			9882 => std_logic_vector(to_unsigned( 215,8)),
			9883 => std_logic_vector(to_unsigned( 168,8)),
			9884 => std_logic_vector(to_unsigned( 79,8)),
			9885 => std_logic_vector(to_unsigned( 232,8)),
			9886 => std_logic_vector(to_unsigned( 133,8)),
			9887 => std_logic_vector(to_unsigned( 153,8)),
			9888 => std_logic_vector(to_unsigned( 198,8)),
			9889 => std_logic_vector(to_unsigned( 140,8)),
			9890 => std_logic_vector(to_unsigned( 219,8)),
			9891 => std_logic_vector(to_unsigned( 50,8)),
			9892 => std_logic_vector(to_unsigned( 238,8)),
			9893 => std_logic_vector(to_unsigned( 79,8)),
			9894 => std_logic_vector(to_unsigned( 141,8)),
			9895 => std_logic_vector(to_unsigned( 78,8)),
			9896 => std_logic_vector(to_unsigned( 191,8)),
			9897 => std_logic_vector(to_unsigned( 11,8)),
			9898 => std_logic_vector(to_unsigned( 199,8)),
			9899 => std_logic_vector(to_unsigned( 183,8)),
			9900 => std_logic_vector(to_unsigned( 225,8)),
			9901 => std_logic_vector(to_unsigned( 116,8)),
			9902 => std_logic_vector(to_unsigned( 15,8)),
			9903 => std_logic_vector(to_unsigned( 224,8)),
			9904 => std_logic_vector(to_unsigned( 137,8)),
			9905 => std_logic_vector(to_unsigned( 237,8)),
			9906 => std_logic_vector(to_unsigned( 37,8)),
			9907 => std_logic_vector(to_unsigned( 172,8)),
			9908 => std_logic_vector(to_unsigned( 108,8)),
			9909 => std_logic_vector(to_unsigned( 73,8)),
			9910 => std_logic_vector(to_unsigned( 160,8)),
			9911 => std_logic_vector(to_unsigned( 195,8)),
			9912 => std_logic_vector(to_unsigned( 113,8)),
			9913 => std_logic_vector(to_unsigned( 183,8)),
			9914 => std_logic_vector(to_unsigned( 116,8)),
			9915 => std_logic_vector(to_unsigned( 55,8)),
			9916 => std_logic_vector(to_unsigned( 102,8)),
			9917 => std_logic_vector(to_unsigned( 168,8)),
			9918 => std_logic_vector(to_unsigned( 195,8)),
			9919 => std_logic_vector(to_unsigned( 61,8)),
			9920 => std_logic_vector(to_unsigned( 221,8)),
			9921 => std_logic_vector(to_unsigned( 146,8)),
			9922 => std_logic_vector(to_unsigned( 33,8)),
			9923 => std_logic_vector(to_unsigned( 72,8)),
			9924 => std_logic_vector(to_unsigned( 117,8)),
			9925 => std_logic_vector(to_unsigned( 28,8)),
			9926 => std_logic_vector(to_unsigned( 195,8)),
			9927 => std_logic_vector(to_unsigned( 234,8)),
			9928 => std_logic_vector(to_unsigned( 191,8)),
			9929 => std_logic_vector(to_unsigned( 14,8)),
			9930 => std_logic_vector(to_unsigned( 158,8)),
			9931 => std_logic_vector(to_unsigned( 173,8)),
			9932 => std_logic_vector(to_unsigned( 142,8)),
			9933 => std_logic_vector(to_unsigned( 123,8)),
			9934 => std_logic_vector(to_unsigned( 142,8)),
			9935 => std_logic_vector(to_unsigned( 64,8)),
			9936 => std_logic_vector(to_unsigned( 153,8)),
			9937 => std_logic_vector(to_unsigned( 168,8)),
			9938 => std_logic_vector(to_unsigned( 161,8)),
			9939 => std_logic_vector(to_unsigned( 106,8)),
			9940 => std_logic_vector(to_unsigned( 82,8)),
			9941 => std_logic_vector(to_unsigned( 72,8)),
			9942 => std_logic_vector(to_unsigned( 221,8)),
			9943 => std_logic_vector(to_unsigned( 29,8)),
			9944 => std_logic_vector(to_unsigned( 58,8)),
			9945 => std_logic_vector(to_unsigned( 16,8)),
			9946 => std_logic_vector(to_unsigned( 91,8)),
			9947 => std_logic_vector(to_unsigned( 26,8)),
			9948 => std_logic_vector(to_unsigned( 158,8)),
			9949 => std_logic_vector(to_unsigned( 10,8)),
			9950 => std_logic_vector(to_unsigned( 24,8)),
			9951 => std_logic_vector(to_unsigned( 128,8)),
			9952 => std_logic_vector(to_unsigned( 23,8)),
			9953 => std_logic_vector(to_unsigned( 242,8)),
			9954 => std_logic_vector(to_unsigned( 33,8)),
			9955 => std_logic_vector(to_unsigned( 247,8)),
			9956 => std_logic_vector(to_unsigned( 221,8)),
			9957 => std_logic_vector(to_unsigned( 195,8)),
			9958 => std_logic_vector(to_unsigned( 191,8)),
			9959 => std_logic_vector(to_unsigned( 96,8)),
			9960 => std_logic_vector(to_unsigned( 207,8)),
			9961 => std_logic_vector(to_unsigned( 71,8)),
			9962 => std_logic_vector(to_unsigned( 109,8)),
			9963 => std_logic_vector(to_unsigned( 77,8)),
			9964 => std_logic_vector(to_unsigned( 165,8)),
			9965 => std_logic_vector(to_unsigned( 33,8)),
			9966 => std_logic_vector(to_unsigned( 89,8)),
			9967 => std_logic_vector(to_unsigned( 218,8)),
			9968 => std_logic_vector(to_unsigned( 173,8)),
			9969 => std_logic_vector(to_unsigned( 142,8)),
			9970 => std_logic_vector(to_unsigned( 254,8)),
			9971 => std_logic_vector(to_unsigned( 157,8)),
			9972 => std_logic_vector(to_unsigned( 114,8)),
			9973 => std_logic_vector(to_unsigned( 108,8)),
			9974 => std_logic_vector(to_unsigned( 62,8)),
			9975 => std_logic_vector(to_unsigned( 121,8)),
			9976 => std_logic_vector(to_unsigned( 128,8)),
			9977 => std_logic_vector(to_unsigned( 178,8)),
			9978 => std_logic_vector(to_unsigned( 217,8)),
			9979 => std_logic_vector(to_unsigned( 95,8)),
			9980 => std_logic_vector(to_unsigned( 4,8)),
			9981 => std_logic_vector(to_unsigned( 240,8)),
			9982 => std_logic_vector(to_unsigned( 220,8)),
			9983 => std_logic_vector(to_unsigned( 177,8)),
			9984 => std_logic_vector(to_unsigned( 27,8)),
			9985 => std_logic_vector(to_unsigned( 109,8)),
			9986 => std_logic_vector(to_unsigned( 138,8)),
			9987 => std_logic_vector(to_unsigned( 81,8)),
			9988 => std_logic_vector(to_unsigned( 138,8)),
			9989 => std_logic_vector(to_unsigned( 102,8)),
			9990 => std_logic_vector(to_unsigned( 39,8)),
			9991 => std_logic_vector(to_unsigned( 90,8)),
			9992 => std_logic_vector(to_unsigned( 41,8)),
			9993 => std_logic_vector(to_unsigned( 60,8)),
			9994 => std_logic_vector(to_unsigned( 8,8)),
			9995 => std_logic_vector(to_unsigned( 128,8)),
			9996 => std_logic_vector(to_unsigned( 43,8)),
			9997 => std_logic_vector(to_unsigned( 131,8)),
			9998 => std_logic_vector(to_unsigned( 79,8)),
			9999 => std_logic_vector(to_unsigned( 143,8)),
			10000 => std_logic_vector(to_unsigned( 168,8)),
			10001 => std_logic_vector(to_unsigned( 2,8)),
			10002 => std_logic_vector(to_unsigned( 205,8)),
			10003 => std_logic_vector(to_unsigned( 51,8)),
			10004 => std_logic_vector(to_unsigned( 221,8)),
			10005 => std_logic_vector(to_unsigned( 135,8)),
			10006 => std_logic_vector(to_unsigned( 124,8)),
			10007 => std_logic_vector(to_unsigned( 123,8)),
			10008 => std_logic_vector(to_unsigned( 7,8)),
			10009 => std_logic_vector(to_unsigned( 134,8)),
			10010 => std_logic_vector(to_unsigned( 154,8)),
			10011 => std_logic_vector(to_unsigned( 166,8)),
			10012 => std_logic_vector(to_unsigned( 62,8)),
			10013 => std_logic_vector(to_unsigned( 184,8)),
			10014 => std_logic_vector(to_unsigned( 209,8)),
			10015 => std_logic_vector(to_unsigned( 228,8)),
			10016 => std_logic_vector(to_unsigned( 25,8)),
			10017 => std_logic_vector(to_unsigned( 231,8)),
			10018 => std_logic_vector(to_unsigned( 135,8)),
			10019 => std_logic_vector(to_unsigned( 3,8)),
			10020 => std_logic_vector(to_unsigned( 199,8)),
			10021 => std_logic_vector(to_unsigned( 220,8)),
			10022 => std_logic_vector(to_unsigned( 141,8)),
			10023 => std_logic_vector(to_unsigned( 121,8)),
			10024 => std_logic_vector(to_unsigned( 114,8)),
			10025 => std_logic_vector(to_unsigned( 170,8)),
			10026 => std_logic_vector(to_unsigned( 232,8)),
			10027 => std_logic_vector(to_unsigned( 45,8)),
			10028 => std_logic_vector(to_unsigned( 63,8)),
			10029 => std_logic_vector(to_unsigned( 147,8)),
			10030 => std_logic_vector(to_unsigned( 189,8)),
			10031 => std_logic_vector(to_unsigned( 179,8)),
			10032 => std_logic_vector(to_unsigned( 211,8)),
			10033 => std_logic_vector(to_unsigned( 28,8)),
			10034 => std_logic_vector(to_unsigned( 47,8)),
			10035 => std_logic_vector(to_unsigned( 23,8)),
			10036 => std_logic_vector(to_unsigned( 220,8)),
			10037 => std_logic_vector(to_unsigned( 9,8)),
			10038 => std_logic_vector(to_unsigned( 178,8)),
			10039 => std_logic_vector(to_unsigned( 253,8)),
			10040 => std_logic_vector(to_unsigned( 78,8)),
			10041 => std_logic_vector(to_unsigned( 254,8)),
			10042 => std_logic_vector(to_unsigned( 154,8)),
			10043 => std_logic_vector(to_unsigned( 169,8)),
			10044 => std_logic_vector(to_unsigned( 147,8)),
			10045 => std_logic_vector(to_unsigned( 128,8)),
			10046 => std_logic_vector(to_unsigned( 62,8)),
			10047 => std_logic_vector(to_unsigned( 197,8)),
			10048 => std_logic_vector(to_unsigned( 4,8)),
			10049 => std_logic_vector(to_unsigned( 48,8)),
			10050 => std_logic_vector(to_unsigned( 73,8)),
			10051 => std_logic_vector(to_unsigned( 167,8)),
			10052 => std_logic_vector(to_unsigned( 56,8)),
			10053 => std_logic_vector(to_unsigned( 34,8)),
			10054 => std_logic_vector(to_unsigned( 212,8)),
			10055 => std_logic_vector(to_unsigned( 53,8)),
			10056 => std_logic_vector(to_unsigned( 214,8)),
			10057 => std_logic_vector(to_unsigned( 155,8)),
			10058 => std_logic_vector(to_unsigned( 108,8)),
			10059 => std_logic_vector(to_unsigned( 150,8)),
			10060 => std_logic_vector(to_unsigned( 57,8)),
			10061 => std_logic_vector(to_unsigned( 60,8)),
			10062 => std_logic_vector(to_unsigned( 53,8)),
			10063 => std_logic_vector(to_unsigned( 163,8)),
			10064 => std_logic_vector(to_unsigned( 57,8)),
			10065 => std_logic_vector(to_unsigned( 82,8)),
			10066 => std_logic_vector(to_unsigned( 198,8)),
			10067 => std_logic_vector(to_unsigned( 246,8)),
			10068 => std_logic_vector(to_unsigned( 100,8)),
			10069 => std_logic_vector(to_unsigned( 49,8)),
			10070 => std_logic_vector(to_unsigned( 105,8)),
			10071 => std_logic_vector(to_unsigned( 92,8)),
			10072 => std_logic_vector(to_unsigned( 44,8)),
			10073 => std_logic_vector(to_unsigned( 240,8)),
			10074 => std_logic_vector(to_unsigned( 250,8)),
			10075 => std_logic_vector(to_unsigned( 144,8)),
			10076 => std_logic_vector(to_unsigned( 198,8)),
			10077 => std_logic_vector(to_unsigned( 248,8)),
			10078 => std_logic_vector(to_unsigned( 4,8)),
			10079 => std_logic_vector(to_unsigned( 174,8)),
			10080 => std_logic_vector(to_unsigned( 30,8)),
			10081 => std_logic_vector(to_unsigned( 178,8)),
			10082 => std_logic_vector(to_unsigned( 250,8)),
			10083 => std_logic_vector(to_unsigned( 254,8)),
			10084 => std_logic_vector(to_unsigned( 67,8)),
			10085 => std_logic_vector(to_unsigned( 218,8)),
			10086 => std_logic_vector(to_unsigned( 86,8)),
			10087 => std_logic_vector(to_unsigned( 105,8)),
			10088 => std_logic_vector(to_unsigned( 135,8)),
			10089 => std_logic_vector(to_unsigned( 182,8)),
			10090 => std_logic_vector(to_unsigned( 151,8)),
			10091 => std_logic_vector(to_unsigned( 69,8)),
			10092 => std_logic_vector(to_unsigned( 64,8)),
			10093 => std_logic_vector(to_unsigned( 203,8)),
			10094 => std_logic_vector(to_unsigned( 246,8)),
			10095 => std_logic_vector(to_unsigned( 84,8)),
			10096 => std_logic_vector(to_unsigned( 248,8)),
			10097 => std_logic_vector(to_unsigned( 98,8)),
			10098 => std_logic_vector(to_unsigned( 2,8)),
			10099 => std_logic_vector(to_unsigned( 172,8)),
			10100 => std_logic_vector(to_unsigned( 127,8)),
			10101 => std_logic_vector(to_unsigned( 139,8)),
			10102 => std_logic_vector(to_unsigned( 203,8)),
			10103 => std_logic_vector(to_unsigned( 12,8)),
			10104 => std_logic_vector(to_unsigned( 255,8)),
			10105 => std_logic_vector(to_unsigned( 5,8)),
			10106 => std_logic_vector(to_unsigned( 154,8)),
			10107 => std_logic_vector(to_unsigned( 233,8)),
			10108 => std_logic_vector(to_unsigned( 253,8)),
			10109 => std_logic_vector(to_unsigned( 247,8)),
			10110 => std_logic_vector(to_unsigned( 52,8)),
			10111 => std_logic_vector(to_unsigned( 132,8)),
			10112 => std_logic_vector(to_unsigned( 222,8)),
			10113 => std_logic_vector(to_unsigned( 92,8)),
			10114 => std_logic_vector(to_unsigned( 14,8)),
			10115 => std_logic_vector(to_unsigned( 109,8)),
			10116 => std_logic_vector(to_unsigned( 154,8)),
			10117 => std_logic_vector(to_unsigned( 236,8)),
			10118 => std_logic_vector(to_unsigned( 102,8)),
			10119 => std_logic_vector(to_unsigned( 199,8)),
			10120 => std_logic_vector(to_unsigned( 50,8)),
			10121 => std_logic_vector(to_unsigned( 51,8)),
			10122 => std_logic_vector(to_unsigned( 22,8)),
			10123 => std_logic_vector(to_unsigned( 57,8)),
			10124 => std_logic_vector(to_unsigned( 213,8)),
			10125 => std_logic_vector(to_unsigned( 117,8)),
			10126 => std_logic_vector(to_unsigned( 31,8)),
			10127 => std_logic_vector(to_unsigned( 0,8)),
			10128 => std_logic_vector(to_unsigned( 129,8)),
			10129 => std_logic_vector(to_unsigned( 200,8)),
			10130 => std_logic_vector(to_unsigned( 46,8)),
			10131 => std_logic_vector(to_unsigned( 132,8)),
			10132 => std_logic_vector(to_unsigned( 232,8)),
			10133 => std_logic_vector(to_unsigned( 226,8)),
			10134 => std_logic_vector(to_unsigned( 23,8)),
			10135 => std_logic_vector(to_unsigned( 83,8)),
			10136 => std_logic_vector(to_unsigned( 56,8)),
			10137 => std_logic_vector(to_unsigned( 203,8)),
			10138 => std_logic_vector(to_unsigned( 125,8)),
			10139 => std_logic_vector(to_unsigned( 8,8)),
			10140 => std_logic_vector(to_unsigned( 127,8)),
			10141 => std_logic_vector(to_unsigned( 156,8)),
			10142 => std_logic_vector(to_unsigned( 127,8)),
			10143 => std_logic_vector(to_unsigned( 0,8)),
			10144 => std_logic_vector(to_unsigned( 212,8)),
			10145 => std_logic_vector(to_unsigned( 36,8)),
			10146 => std_logic_vector(to_unsigned( 196,8)),
			10147 => std_logic_vector(to_unsigned( 204,8)),
			10148 => std_logic_vector(to_unsigned( 246,8)),
			10149 => std_logic_vector(to_unsigned( 6,8)),
			10150 => std_logic_vector(to_unsigned( 242,8)),
			10151 => std_logic_vector(to_unsigned( 151,8)),
			10152 => std_logic_vector(to_unsigned( 104,8)),
			10153 => std_logic_vector(to_unsigned( 71,8)),
			10154 => std_logic_vector(to_unsigned( 18,8)),
			10155 => std_logic_vector(to_unsigned( 176,8)),
			10156 => std_logic_vector(to_unsigned( 21,8)),
			10157 => std_logic_vector(to_unsigned( 233,8)),
			10158 => std_logic_vector(to_unsigned( 179,8)),
			10159 => std_logic_vector(to_unsigned( 73,8)),
			10160 => std_logic_vector(to_unsigned( 204,8)),
			10161 => std_logic_vector(to_unsigned( 132,8)),
			10162 => std_logic_vector(to_unsigned( 67,8)),
			10163 => std_logic_vector(to_unsigned( 232,8)),
			10164 => std_logic_vector(to_unsigned( 222,8)),
			10165 => std_logic_vector(to_unsigned( 6,8)),
			10166 => std_logic_vector(to_unsigned( 81,8)),
			10167 => std_logic_vector(to_unsigned( 118,8)),
			10168 => std_logic_vector(to_unsigned( 203,8)),
			10169 => std_logic_vector(to_unsigned( 18,8)),
			10170 => std_logic_vector(to_unsigned( 244,8)),
			10171 => std_logic_vector(to_unsigned( 188,8)),
			10172 => std_logic_vector(to_unsigned( 75,8)),
			10173 => std_logic_vector(to_unsigned( 53,8)),
			10174 => std_logic_vector(to_unsigned( 208,8)),
			10175 => std_logic_vector(to_unsigned( 36,8)),
			10176 => std_logic_vector(to_unsigned( 36,8)),
			10177 => std_logic_vector(to_unsigned( 114,8)),
			10178 => std_logic_vector(to_unsigned( 247,8)),
			10179 => std_logic_vector(to_unsigned( 128,8)),
			10180 => std_logic_vector(to_unsigned( 230,8)),
			10181 => std_logic_vector(to_unsigned( 159,8)),
			10182 => std_logic_vector(to_unsigned( 159,8)),
			10183 => std_logic_vector(to_unsigned( 84,8)),
			10184 => std_logic_vector(to_unsigned( 208,8)),
			10185 => std_logic_vector(to_unsigned( 204,8)),
			10186 => std_logic_vector(to_unsigned( 87,8)),
			10187 => std_logic_vector(to_unsigned( 223,8)),
			10188 => std_logic_vector(to_unsigned( 161,8)),
			10189 => std_logic_vector(to_unsigned( 114,8)),
			10190 => std_logic_vector(to_unsigned( 187,8)),
			10191 => std_logic_vector(to_unsigned( 110,8)),
			10192 => std_logic_vector(to_unsigned( 252,8)),
			10193 => std_logic_vector(to_unsigned( 162,8)),
			10194 => std_logic_vector(to_unsigned( 244,8)),
			10195 => std_logic_vector(to_unsigned( 2,8)),
			10196 => std_logic_vector(to_unsigned( 156,8)),
			10197 => std_logic_vector(to_unsigned( 253,8)),
			10198 => std_logic_vector(to_unsigned( 108,8)),
			10199 => std_logic_vector(to_unsigned( 148,8)),
			10200 => std_logic_vector(to_unsigned( 198,8)),
			10201 => std_logic_vector(to_unsigned( 143,8)),
			10202 => std_logic_vector(to_unsigned( 40,8)),
			10203 => std_logic_vector(to_unsigned( 201,8)),
			10204 => std_logic_vector(to_unsigned( 198,8)),
			10205 => std_logic_vector(to_unsigned( 98,8)),
			10206 => std_logic_vector(to_unsigned( 134,8)),
			10207 => std_logic_vector(to_unsigned( 218,8)),
			10208 => std_logic_vector(to_unsigned( 229,8)),
			10209 => std_logic_vector(to_unsigned( 5,8)),
			10210 => std_logic_vector(to_unsigned( 82,8)),
			10211 => std_logic_vector(to_unsigned( 226,8)),
			10212 => std_logic_vector(to_unsigned( 102,8)),
			10213 => std_logic_vector(to_unsigned( 181,8)),
			10214 => std_logic_vector(to_unsigned( 190,8)),
			10215 => std_logic_vector(to_unsigned( 77,8)),
			10216 => std_logic_vector(to_unsigned( 211,8)),
			10217 => std_logic_vector(to_unsigned( 180,8)),
			10218 => std_logic_vector(to_unsigned( 55,8)),
			10219 => std_logic_vector(to_unsigned( 209,8)),
			10220 => std_logic_vector(to_unsigned( 216,8)),
			10221 => std_logic_vector(to_unsigned( 188,8)),
			10222 => std_logic_vector(to_unsigned( 211,8)),
			10223 => std_logic_vector(to_unsigned( 94,8)),
			10224 => std_logic_vector(to_unsigned( 177,8)),
			10225 => std_logic_vector(to_unsigned( 254,8)),
			10226 => std_logic_vector(to_unsigned( 174,8)),
			10227 => std_logic_vector(to_unsigned( 49,8)),
			10228 => std_logic_vector(to_unsigned( 231,8)),
			10229 => std_logic_vector(to_unsigned( 101,8)),
			10230 => std_logic_vector(to_unsigned( 193,8)),
			10231 => std_logic_vector(to_unsigned( 92,8)),
			10232 => std_logic_vector(to_unsigned( 149,8)),
			10233 => std_logic_vector(to_unsigned( 219,8)),
			10234 => std_logic_vector(to_unsigned( 67,8)),
			10235 => std_logic_vector(to_unsigned( 18,8)),
			10236 => std_logic_vector(to_unsigned( 100,8)),
			10237 => std_logic_vector(to_unsigned( 0,8)),
			10238 => std_logic_vector(to_unsigned( 142,8)),
			10239 => std_logic_vector(to_unsigned( 59,8)),
			10240 => std_logic_vector(to_unsigned( 243,8)),
			10241 => std_logic_vector(to_unsigned( 26,8)),
			10242 => std_logic_vector(to_unsigned( 254,8)),
			10243 => std_logic_vector(to_unsigned( 219,8)),
			10244 => std_logic_vector(to_unsigned( 181,8)),
			10245 => std_logic_vector(to_unsigned( 127,8)),
			10246 => std_logic_vector(to_unsigned( 165,8)),
			10247 => std_logic_vector(to_unsigned( 24,8)),
			10248 => std_logic_vector(to_unsigned( 193,8)),
			10249 => std_logic_vector(to_unsigned( 234,8)),
			10250 => std_logic_vector(to_unsigned( 58,8)),
			10251 => std_logic_vector(to_unsigned( 25,8)),
			10252 => std_logic_vector(to_unsigned( 94,8)),
			10253 => std_logic_vector(to_unsigned( 118,8)),
			10254 => std_logic_vector(to_unsigned( 63,8)),
			10255 => std_logic_vector(to_unsigned( 39,8)),
			10256 => std_logic_vector(to_unsigned( 43,8)),
			10257 => std_logic_vector(to_unsigned( 129,8)),
			10258 => std_logic_vector(to_unsigned( 80,8)),
			10259 => std_logic_vector(to_unsigned( 198,8)),
			10260 => std_logic_vector(to_unsigned( 33,8)),
			10261 => std_logic_vector(to_unsigned( 144,8)),
			10262 => std_logic_vector(to_unsigned( 31,8)),
			10263 => std_logic_vector(to_unsigned( 205,8)),
			10264 => std_logic_vector(to_unsigned( 190,8)),
			10265 => std_logic_vector(to_unsigned( 127,8)),
			10266 => std_logic_vector(to_unsigned( 45,8)),
			10267 => std_logic_vector(to_unsigned( 205,8)),
			10268 => std_logic_vector(to_unsigned( 150,8)),
			10269 => std_logic_vector(to_unsigned( 1,8)),
			10270 => std_logic_vector(to_unsigned( 213,8)),
			10271 => std_logic_vector(to_unsigned( 214,8)),
			10272 => std_logic_vector(to_unsigned( 152,8)),
			10273 => std_logic_vector(to_unsigned( 75,8)),
			10274 => std_logic_vector(to_unsigned( 31,8)),
			10275 => std_logic_vector(to_unsigned( 27,8)),
			10276 => std_logic_vector(to_unsigned( 139,8)),
			10277 => std_logic_vector(to_unsigned( 74,8)),
			10278 => std_logic_vector(to_unsigned( 106,8)),
			10279 => std_logic_vector(to_unsigned( 170,8)),
			10280 => std_logic_vector(to_unsigned( 151,8)),
			10281 => std_logic_vector(to_unsigned( 131,8)),
			10282 => std_logic_vector(to_unsigned( 122,8)),
			10283 => std_logic_vector(to_unsigned( 140,8)),
			10284 => std_logic_vector(to_unsigned( 11,8)),
			10285 => std_logic_vector(to_unsigned( 169,8)),
			10286 => std_logic_vector(to_unsigned( 249,8)),
			10287 => std_logic_vector(to_unsigned( 134,8)),
			10288 => std_logic_vector(to_unsigned( 43,8)),
			10289 => std_logic_vector(to_unsigned( 238,8)),
			10290 => std_logic_vector(to_unsigned( 29,8)),
			10291 => std_logic_vector(to_unsigned( 176,8)),
			10292 => std_logic_vector(to_unsigned( 226,8)),
			10293 => std_logic_vector(to_unsigned( 227,8)),
			10294 => std_logic_vector(to_unsigned( 103,8)),
			10295 => std_logic_vector(to_unsigned( 67,8)),
			10296 => std_logic_vector(to_unsigned( 156,8)),
			10297 => std_logic_vector(to_unsigned( 125,8)),
			10298 => std_logic_vector(to_unsigned( 143,8)),
			10299 => std_logic_vector(to_unsigned( 81,8)),
			10300 => std_logic_vector(to_unsigned( 26,8)),
			10301 => std_logic_vector(to_unsigned( 168,8)),
			10302 => std_logic_vector(to_unsigned( 39,8)),
			10303 => std_logic_vector(to_unsigned( 184,8)),
			10304 => std_logic_vector(to_unsigned( 190,8)),
			10305 => std_logic_vector(to_unsigned( 32,8)),
			10306 => std_logic_vector(to_unsigned( 75,8)),
			10307 => std_logic_vector(to_unsigned( 88,8)),
			10308 => std_logic_vector(to_unsigned( 194,8)),
			10309 => std_logic_vector(to_unsigned( 223,8)),
			10310 => std_logic_vector(to_unsigned( 223,8)),
			10311 => std_logic_vector(to_unsigned( 111,8)),
			10312 => std_logic_vector(to_unsigned( 84,8)),
			10313 => std_logic_vector(to_unsigned( 79,8)),
			10314 => std_logic_vector(to_unsigned( 124,8)),
			10315 => std_logic_vector(to_unsigned( 192,8)),
			10316 => std_logic_vector(to_unsigned( 247,8)),
			10317 => std_logic_vector(to_unsigned( 202,8)),
			10318 => std_logic_vector(to_unsigned( 7,8)),
			10319 => std_logic_vector(to_unsigned( 81,8)),
			10320 => std_logic_vector(to_unsigned( 101,8)),
			10321 => std_logic_vector(to_unsigned( 177,8)),
			10322 => std_logic_vector(to_unsigned( 250,8)),
			10323 => std_logic_vector(to_unsigned( 149,8)),
			10324 => std_logic_vector(to_unsigned( 127,8)),
			10325 => std_logic_vector(to_unsigned( 38,8)),
			10326 => std_logic_vector(to_unsigned( 166,8)),
			10327 => std_logic_vector(to_unsigned( 158,8)),
			10328 => std_logic_vector(to_unsigned( 61,8)),
			10329 => std_logic_vector(to_unsigned( 187,8)),
			10330 => std_logic_vector(to_unsigned( 56,8)),
			10331 => std_logic_vector(to_unsigned( 171,8)),
			10332 => std_logic_vector(to_unsigned( 33,8)),
			10333 => std_logic_vector(to_unsigned( 203,8)),
			10334 => std_logic_vector(to_unsigned( 208,8)),
			10335 => std_logic_vector(to_unsigned( 105,8)),
			10336 => std_logic_vector(to_unsigned( 126,8)),
			10337 => std_logic_vector(to_unsigned( 92,8)),
			10338 => std_logic_vector(to_unsigned( 99,8)),
			10339 => std_logic_vector(to_unsigned( 226,8)),
			10340 => std_logic_vector(to_unsigned( 21,8)),
			10341 => std_logic_vector(to_unsigned( 59,8)),
			10342 => std_logic_vector(to_unsigned( 250,8)),
			10343 => std_logic_vector(to_unsigned( 210,8)),
			10344 => std_logic_vector(to_unsigned( 208,8)),
			10345 => std_logic_vector(to_unsigned( 231,8)),
			10346 => std_logic_vector(to_unsigned( 122,8)),
			10347 => std_logic_vector(to_unsigned( 51,8)),
			10348 => std_logic_vector(to_unsigned( 47,8)),
			10349 => std_logic_vector(to_unsigned( 226,8)),
			10350 => std_logic_vector(to_unsigned( 72,8)),
			10351 => std_logic_vector(to_unsigned( 43,8)),
			10352 => std_logic_vector(to_unsigned( 252,8)),
			10353 => std_logic_vector(to_unsigned( 161,8)),
			10354 => std_logic_vector(to_unsigned( 123,8)),
			10355 => std_logic_vector(to_unsigned( 242,8)),
			10356 => std_logic_vector(to_unsigned( 83,8)),
			10357 => std_logic_vector(to_unsigned( 20,8)),
			10358 => std_logic_vector(to_unsigned( 46,8)),
			10359 => std_logic_vector(to_unsigned( 0,8)),
			10360 => std_logic_vector(to_unsigned( 38,8)),
			10361 => std_logic_vector(to_unsigned( 35,8)),
			10362 => std_logic_vector(to_unsigned( 111,8)),
			10363 => std_logic_vector(to_unsigned( 74,8)),
			10364 => std_logic_vector(to_unsigned( 218,8)),
			10365 => std_logic_vector(to_unsigned( 195,8)),
			10366 => std_logic_vector(to_unsigned( 36,8)),
			10367 => std_logic_vector(to_unsigned( 111,8)),
			10368 => std_logic_vector(to_unsigned( 199,8)),
			10369 => std_logic_vector(to_unsigned( 137,8)),
			10370 => std_logic_vector(to_unsigned( 194,8)),
			10371 => std_logic_vector(to_unsigned( 42,8)),
			10372 => std_logic_vector(to_unsigned( 4,8)),
			10373 => std_logic_vector(to_unsigned( 76,8)),
			10374 => std_logic_vector(to_unsigned( 147,8)),
			10375 => std_logic_vector(to_unsigned( 245,8)),
			10376 => std_logic_vector(to_unsigned( 33,8)),
			10377 => std_logic_vector(to_unsigned( 118,8)),
			10378 => std_logic_vector(to_unsigned( 99,8)),
			10379 => std_logic_vector(to_unsigned( 84,8)),
			10380 => std_logic_vector(to_unsigned( 91,8)),
			10381 => std_logic_vector(to_unsigned( 84,8)),
			10382 => std_logic_vector(to_unsigned( 109,8)),
			10383 => std_logic_vector(to_unsigned( 112,8)),
			10384 => std_logic_vector(to_unsigned( 43,8)),
			10385 => std_logic_vector(to_unsigned( 77,8)),
			10386 => std_logic_vector(to_unsigned( 56,8)),
			10387 => std_logic_vector(to_unsigned( 153,8)),
			10388 => std_logic_vector(to_unsigned( 228,8)),
			10389 => std_logic_vector(to_unsigned( 135,8)),
			10390 => std_logic_vector(to_unsigned( 96,8)),
			10391 => std_logic_vector(to_unsigned( 166,8)),
			10392 => std_logic_vector(to_unsigned( 20,8)),
			10393 => std_logic_vector(to_unsigned( 204,8)),
			10394 => std_logic_vector(to_unsigned( 136,8)),
			10395 => std_logic_vector(to_unsigned( 52,8)),
			10396 => std_logic_vector(to_unsigned( 133,8)),
			10397 => std_logic_vector(to_unsigned( 121,8)),
			10398 => std_logic_vector(to_unsigned( 154,8)),
			10399 => std_logic_vector(to_unsigned( 244,8)),
			10400 => std_logic_vector(to_unsigned( 208,8)),
			10401 => std_logic_vector(to_unsigned( 140,8)),
			10402 => std_logic_vector(to_unsigned( 3,8)),
			10403 => std_logic_vector(to_unsigned( 84,8)),
			10404 => std_logic_vector(to_unsigned( 196,8)),
			10405 => std_logic_vector(to_unsigned( 71,8)),
			10406 => std_logic_vector(to_unsigned( 210,8)),
			10407 => std_logic_vector(to_unsigned( 186,8)),
			10408 => std_logic_vector(to_unsigned( 133,8)),
			10409 => std_logic_vector(to_unsigned( 116,8)),
			10410 => std_logic_vector(to_unsigned( 229,8)),
			10411 => std_logic_vector(to_unsigned( 17,8)),
			10412 => std_logic_vector(to_unsigned( 93,8)),
			10413 => std_logic_vector(to_unsigned( 17,8)),
			10414 => std_logic_vector(to_unsigned( 93,8)),
			10415 => std_logic_vector(to_unsigned( 168,8)),
			10416 => std_logic_vector(to_unsigned( 208,8)),
			10417 => std_logic_vector(to_unsigned( 212,8)),
			10418 => std_logic_vector(to_unsigned( 59,8)),
			10419 => std_logic_vector(to_unsigned( 184,8)),
			10420 => std_logic_vector(to_unsigned( 166,8)),
			10421 => std_logic_vector(to_unsigned( 91,8)),
			10422 => std_logic_vector(to_unsigned( 18,8)),
			10423 => std_logic_vector(to_unsigned( 91,8)),
			10424 => std_logic_vector(to_unsigned( 169,8)),
			10425 => std_logic_vector(to_unsigned( 223,8)),
			10426 => std_logic_vector(to_unsigned( 227,8)),
			10427 => std_logic_vector(to_unsigned( 116,8)),
			10428 => std_logic_vector(to_unsigned( 89,8)),
			10429 => std_logic_vector(to_unsigned( 4,8)),
			10430 => std_logic_vector(to_unsigned( 251,8)),
			10431 => std_logic_vector(to_unsigned( 109,8)),
			10432 => std_logic_vector(to_unsigned( 93,8)),
			10433 => std_logic_vector(to_unsigned( 108,8)),
			10434 => std_logic_vector(to_unsigned( 251,8)),
			10435 => std_logic_vector(to_unsigned( 75,8)),
			10436 => std_logic_vector(to_unsigned( 48,8)),
			10437 => std_logic_vector(to_unsigned( 196,8)),
			10438 => std_logic_vector(to_unsigned( 212,8)),
			10439 => std_logic_vector(to_unsigned( 35,8)),
			10440 => std_logic_vector(to_unsigned( 96,8)),
			10441 => std_logic_vector(to_unsigned( 225,8)),
			10442 => std_logic_vector(to_unsigned( 240,8)),
			10443 => std_logic_vector(to_unsigned( 3,8)),
			10444 => std_logic_vector(to_unsigned( 29,8)),
			10445 => std_logic_vector(to_unsigned( 102,8)),
			10446 => std_logic_vector(to_unsigned( 80,8)),
			10447 => std_logic_vector(to_unsigned( 23,8)),
			10448 => std_logic_vector(to_unsigned( 39,8)),
			10449 => std_logic_vector(to_unsigned( 158,8)),
			10450 => std_logic_vector(to_unsigned( 188,8)),
			10451 => std_logic_vector(to_unsigned( 143,8)),
			10452 => std_logic_vector(to_unsigned( 146,8)),
			10453 => std_logic_vector(to_unsigned( 89,8)),
			10454 => std_logic_vector(to_unsigned( 117,8)),
			10455 => std_logic_vector(to_unsigned( 117,8)),
			10456 => std_logic_vector(to_unsigned( 114,8)),
			10457 => std_logic_vector(to_unsigned( 61,8)),
			10458 => std_logic_vector(to_unsigned( 39,8)),
			10459 => std_logic_vector(to_unsigned( 253,8)),
			10460 => std_logic_vector(to_unsigned( 112,8)),
			10461 => std_logic_vector(to_unsigned( 137,8)),
			10462 => std_logic_vector(to_unsigned( 80,8)),
			10463 => std_logic_vector(to_unsigned( 122,8)),
			10464 => std_logic_vector(to_unsigned( 40,8)),
			10465 => std_logic_vector(to_unsigned( 243,8)),
			10466 => std_logic_vector(to_unsigned( 182,8)),
			10467 => std_logic_vector(to_unsigned( 104,8)),
			10468 => std_logic_vector(to_unsigned( 164,8)),
			10469 => std_logic_vector(to_unsigned( 124,8)),
			10470 => std_logic_vector(to_unsigned( 234,8)),
			10471 => std_logic_vector(to_unsigned( 223,8)),
			10472 => std_logic_vector(to_unsigned( 146,8)),
			10473 => std_logic_vector(to_unsigned( 71,8)),
			10474 => std_logic_vector(to_unsigned( 24,8)),
			10475 => std_logic_vector(to_unsigned( 81,8)),
			10476 => std_logic_vector(to_unsigned( 255,8)),
			10477 => std_logic_vector(to_unsigned( 254,8)),
			10478 => std_logic_vector(to_unsigned( 146,8)),
			10479 => std_logic_vector(to_unsigned( 87,8)),
			10480 => std_logic_vector(to_unsigned( 107,8)),
			10481 => std_logic_vector(to_unsigned( 207,8)),
			10482 => std_logic_vector(to_unsigned( 35,8)),
			10483 => std_logic_vector(to_unsigned( 216,8)),
			10484 => std_logic_vector(to_unsigned( 121,8)),
			10485 => std_logic_vector(to_unsigned( 114,8)),
			10486 => std_logic_vector(to_unsigned( 222,8)),
			10487 => std_logic_vector(to_unsigned( 235,8)),
			10488 => std_logic_vector(to_unsigned( 236,8)),
			10489 => std_logic_vector(to_unsigned( 65,8)),
			10490 => std_logic_vector(to_unsigned( 86,8)),
			10491 => std_logic_vector(to_unsigned( 57,8)),
			10492 => std_logic_vector(to_unsigned( 103,8)),
			10493 => std_logic_vector(to_unsigned( 102,8)),
			10494 => std_logic_vector(to_unsigned( 207,8)),
			10495 => std_logic_vector(to_unsigned( 56,8)),
			10496 => std_logic_vector(to_unsigned( 66,8)),
			10497 => std_logic_vector(to_unsigned( 139,8)),
			10498 => std_logic_vector(to_unsigned( 25,8)),
			10499 => std_logic_vector(to_unsigned( 88,8)),
			10500 => std_logic_vector(to_unsigned( 109,8)),
			10501 => std_logic_vector(to_unsigned( 16,8)),
			10502 => std_logic_vector(to_unsigned( 197,8)),
			10503 => std_logic_vector(to_unsigned( 224,8)),
			10504 => std_logic_vector(to_unsigned( 152,8)),
			10505 => std_logic_vector(to_unsigned( 97,8)),
			10506 => std_logic_vector(to_unsigned( 34,8)),
			10507 => std_logic_vector(to_unsigned( 47,8)),
			10508 => std_logic_vector(to_unsigned( 112,8)),
			10509 => std_logic_vector(to_unsigned( 86,8)),
			10510 => std_logic_vector(to_unsigned( 215,8)),
			10511 => std_logic_vector(to_unsigned( 211,8)),
			10512 => std_logic_vector(to_unsigned( 72,8)),
			10513 => std_logic_vector(to_unsigned( 57,8)),
			10514 => std_logic_vector(to_unsigned( 64,8)),
			10515 => std_logic_vector(to_unsigned( 143,8)),
			10516 => std_logic_vector(to_unsigned( 95,8)),
			10517 => std_logic_vector(to_unsigned( 37,8)),
			10518 => std_logic_vector(to_unsigned( 254,8)),
			10519 => std_logic_vector(to_unsigned( 100,8)),
			10520 => std_logic_vector(to_unsigned( 209,8)),
			10521 => std_logic_vector(to_unsigned( 249,8)),
			10522 => std_logic_vector(to_unsigned( 178,8)),
			10523 => std_logic_vector(to_unsigned( 75,8)),
			10524 => std_logic_vector(to_unsigned( 147,8)),
			10525 => std_logic_vector(to_unsigned( 104,8)),
			10526 => std_logic_vector(to_unsigned( 166,8)),
			10527 => std_logic_vector(to_unsigned( 250,8)),
			10528 => std_logic_vector(to_unsigned( 216,8)),
			10529 => std_logic_vector(to_unsigned( 49,8)),
			10530 => std_logic_vector(to_unsigned( 193,8)),
			10531 => std_logic_vector(to_unsigned( 52,8)),
			10532 => std_logic_vector(to_unsigned( 150,8)),
			10533 => std_logic_vector(to_unsigned( 13,8)),
			10534 => std_logic_vector(to_unsigned( 75,8)),
			10535 => std_logic_vector(to_unsigned( 31,8)),
			10536 => std_logic_vector(to_unsigned( 247,8)),
			10537 => std_logic_vector(to_unsigned( 152,8)),
			10538 => std_logic_vector(to_unsigned( 201,8)),
			10539 => std_logic_vector(to_unsigned( 38,8)),
			10540 => std_logic_vector(to_unsigned( 128,8)),
			10541 => std_logic_vector(to_unsigned( 203,8)),
			10542 => std_logic_vector(to_unsigned( 136,8)),
			10543 => std_logic_vector(to_unsigned( 141,8)),
			10544 => std_logic_vector(to_unsigned( 72,8)),
			10545 => std_logic_vector(to_unsigned( 13,8)),
			10546 => std_logic_vector(to_unsigned( 186,8)),
			10547 => std_logic_vector(to_unsigned( 67,8)),
			10548 => std_logic_vector(to_unsigned( 158,8)),
			10549 => std_logic_vector(to_unsigned( 139,8)),
			10550 => std_logic_vector(to_unsigned( 168,8)),
			10551 => std_logic_vector(to_unsigned( 229,8)),
			10552 => std_logic_vector(to_unsigned( 96,8)),
			10553 => std_logic_vector(to_unsigned( 169,8)),
			10554 => std_logic_vector(to_unsigned( 171,8)),
			10555 => std_logic_vector(to_unsigned( 50,8)),
			10556 => std_logic_vector(to_unsigned( 42,8)),
			10557 => std_logic_vector(to_unsigned( 145,8)),
			10558 => std_logic_vector(to_unsigned( 1,8)),
			10559 => std_logic_vector(to_unsigned( 164,8)),
			10560 => std_logic_vector(to_unsigned( 96,8)),
			10561 => std_logic_vector(to_unsigned( 179,8)),
			10562 => std_logic_vector(to_unsigned( 86,8)),
			10563 => std_logic_vector(to_unsigned( 14,8)),
			10564 => std_logic_vector(to_unsigned( 62,8)),
			10565 => std_logic_vector(to_unsigned( 16,8)),
			10566 => std_logic_vector(to_unsigned( 92,8)),
			10567 => std_logic_vector(to_unsigned( 175,8)),
			10568 => std_logic_vector(to_unsigned( 84,8)),
			10569 => std_logic_vector(to_unsigned( 153,8)),
			10570 => std_logic_vector(to_unsigned( 4,8)),
			10571 => std_logic_vector(to_unsigned( 131,8)),
			10572 => std_logic_vector(to_unsigned( 72,8)),
			10573 => std_logic_vector(to_unsigned( 203,8)),
			10574 => std_logic_vector(to_unsigned( 8,8)),
			10575 => std_logic_vector(to_unsigned( 111,8)),
			10576 => std_logic_vector(to_unsigned( 251,8)),
			10577 => std_logic_vector(to_unsigned( 214,8)),
			10578 => std_logic_vector(to_unsigned( 16,8)),
			10579 => std_logic_vector(to_unsigned( 233,8)),
			10580 => std_logic_vector(to_unsigned( 24,8)),
			10581 => std_logic_vector(to_unsigned( 53,8)),
			10582 => std_logic_vector(to_unsigned( 215,8)),
			10583 => std_logic_vector(to_unsigned( 153,8)),
			10584 => std_logic_vector(to_unsigned( 186,8)),
			10585 => std_logic_vector(to_unsigned( 96,8)),
			10586 => std_logic_vector(to_unsigned( 31,8)),
			10587 => std_logic_vector(to_unsigned( 207,8)),
			10588 => std_logic_vector(to_unsigned( 117,8)),
			10589 => std_logic_vector(to_unsigned( 2,8)),
			10590 => std_logic_vector(to_unsigned( 254,8)),
			10591 => std_logic_vector(to_unsigned( 100,8)),
			10592 => std_logic_vector(to_unsigned( 136,8)),
			10593 => std_logic_vector(to_unsigned( 6,8)),
			10594 => std_logic_vector(to_unsigned( 39,8)),
			10595 => std_logic_vector(to_unsigned( 111,8)),
			10596 => std_logic_vector(to_unsigned( 156,8)),
			10597 => std_logic_vector(to_unsigned( 240,8)),
			10598 => std_logic_vector(to_unsigned( 113,8)),
			10599 => std_logic_vector(to_unsigned( 165,8)),
			10600 => std_logic_vector(to_unsigned( 156,8)),
			10601 => std_logic_vector(to_unsigned( 165,8)),
			10602 => std_logic_vector(to_unsigned( 59,8)),
			10603 => std_logic_vector(to_unsigned( 72,8)),
			10604 => std_logic_vector(to_unsigned( 112,8)),
			10605 => std_logic_vector(to_unsigned( 93,8)),
			10606 => std_logic_vector(to_unsigned( 226,8)),
			10607 => std_logic_vector(to_unsigned( 130,8)),
			10608 => std_logic_vector(to_unsigned( 232,8)),
			10609 => std_logic_vector(to_unsigned( 73,8)),
			10610 => std_logic_vector(to_unsigned( 34,8)),
			10611 => std_logic_vector(to_unsigned( 139,8)),
			10612 => std_logic_vector(to_unsigned( 205,8)),
			10613 => std_logic_vector(to_unsigned( 218,8)),
			10614 => std_logic_vector(to_unsigned( 95,8)),
			10615 => std_logic_vector(to_unsigned( 242,8)),
			10616 => std_logic_vector(to_unsigned( 209,8)),
			10617 => std_logic_vector(to_unsigned( 216,8)),
			10618 => std_logic_vector(to_unsigned( 25,8)),
			10619 => std_logic_vector(to_unsigned( 107,8)),
			10620 => std_logic_vector(to_unsigned( 239,8)),
			10621 => std_logic_vector(to_unsigned( 86,8)),
			10622 => std_logic_vector(to_unsigned( 230,8)),
			10623 => std_logic_vector(to_unsigned( 119,8)),
			10624 => std_logic_vector(to_unsigned( 17,8)),
			10625 => std_logic_vector(to_unsigned( 207,8)),
			10626 => std_logic_vector(to_unsigned( 4,8)),
			10627 => std_logic_vector(to_unsigned( 222,8)),
			10628 => std_logic_vector(to_unsigned( 18,8)),
			10629 => std_logic_vector(to_unsigned( 137,8)),
			10630 => std_logic_vector(to_unsigned( 61,8)),
			10631 => std_logic_vector(to_unsigned( 100,8)),
			10632 => std_logic_vector(to_unsigned( 30,8)),
			10633 => std_logic_vector(to_unsigned( 187,8)),
			10634 => std_logic_vector(to_unsigned( 67,8)),
			10635 => std_logic_vector(to_unsigned( 175,8)),
			10636 => std_logic_vector(to_unsigned( 150,8)),
			10637 => std_logic_vector(to_unsigned( 90,8)),
			10638 => std_logic_vector(to_unsigned( 154,8)),
			10639 => std_logic_vector(to_unsigned( 14,8)),
			10640 => std_logic_vector(to_unsigned( 71,8)),
			10641 => std_logic_vector(to_unsigned( 234,8)),
			10642 => std_logic_vector(to_unsigned( 165,8)),
			10643 => std_logic_vector(to_unsigned( 215,8)),
			10644 => std_logic_vector(to_unsigned( 21,8)),
			10645 => std_logic_vector(to_unsigned( 38,8)),
			10646 => std_logic_vector(to_unsigned( 175,8)),
			10647 => std_logic_vector(to_unsigned( 237,8)),
			10648 => std_logic_vector(to_unsigned( 71,8)),
			10649 => std_logic_vector(to_unsigned( 36,8)),
			10650 => std_logic_vector(to_unsigned( 45,8)),
			10651 => std_logic_vector(to_unsigned( 80,8)),
			10652 => std_logic_vector(to_unsigned( 52,8)),
			10653 => std_logic_vector(to_unsigned( 24,8)),
			10654 => std_logic_vector(to_unsigned( 3,8)),
			10655 => std_logic_vector(to_unsigned( 40,8)),
			10656 => std_logic_vector(to_unsigned( 203,8)),
			10657 => std_logic_vector(to_unsigned( 23,8)),
			10658 => std_logic_vector(to_unsigned( 197,8)),
			10659 => std_logic_vector(to_unsigned( 59,8)),
			10660 => std_logic_vector(to_unsigned( 66,8)),
			10661 => std_logic_vector(to_unsigned( 158,8)),
			10662 => std_logic_vector(to_unsigned( 41,8)),
			10663 => std_logic_vector(to_unsigned( 63,8)),
			10664 => std_logic_vector(to_unsigned( 212,8)),
			10665 => std_logic_vector(to_unsigned( 224,8)),
			10666 => std_logic_vector(to_unsigned( 228,8)),
			10667 => std_logic_vector(to_unsigned( 233,8)),
			10668 => std_logic_vector(to_unsigned( 198,8)),
			10669 => std_logic_vector(to_unsigned( 21,8)),
			10670 => std_logic_vector(to_unsigned( 131,8)),
			10671 => std_logic_vector(to_unsigned( 111,8)),
			10672 => std_logic_vector(to_unsigned( 51,8)),
			10673 => std_logic_vector(to_unsigned( 249,8)),
			10674 => std_logic_vector(to_unsigned( 44,8)),
			10675 => std_logic_vector(to_unsigned( 239,8)),
			10676 => std_logic_vector(to_unsigned( 74,8)),
			10677 => std_logic_vector(to_unsigned( 235,8)),
			10678 => std_logic_vector(to_unsigned( 156,8)),
			10679 => std_logic_vector(to_unsigned( 113,8)),
			10680 => std_logic_vector(to_unsigned( 120,8)),
			10681 => std_logic_vector(to_unsigned( 109,8)),
			10682 => std_logic_vector(to_unsigned( 187,8)),
			10683 => std_logic_vector(to_unsigned( 28,8)),
			10684 => std_logic_vector(to_unsigned( 166,8)),
			10685 => std_logic_vector(to_unsigned( 87,8)),
			10686 => std_logic_vector(to_unsigned( 96,8)),
			10687 => std_logic_vector(to_unsigned( 221,8)),
			10688 => std_logic_vector(to_unsigned( 191,8)),
			10689 => std_logic_vector(to_unsigned( 103,8)),
			10690 => std_logic_vector(to_unsigned( 4,8)),
			10691 => std_logic_vector(to_unsigned( 24,8)),
			10692 => std_logic_vector(to_unsigned( 52,8)),
			10693 => std_logic_vector(to_unsigned( 27,8)),
			10694 => std_logic_vector(to_unsigned( 212,8)),
			10695 => std_logic_vector(to_unsigned( 111,8)),
			10696 => std_logic_vector(to_unsigned( 36,8)),
			10697 => std_logic_vector(to_unsigned( 162,8)),
			10698 => std_logic_vector(to_unsigned( 91,8)),
			10699 => std_logic_vector(to_unsigned( 163,8)),
			10700 => std_logic_vector(to_unsigned( 194,8)),
			10701 => std_logic_vector(to_unsigned( 150,8)),
			10702 => std_logic_vector(to_unsigned( 24,8)),
			10703 => std_logic_vector(to_unsigned( 156,8)),
			10704 => std_logic_vector(to_unsigned( 176,8)),
			10705 => std_logic_vector(to_unsigned( 10,8)),
			10706 => std_logic_vector(to_unsigned( 175,8)),
			10707 => std_logic_vector(to_unsigned( 224,8)),
			10708 => std_logic_vector(to_unsigned( 169,8)),
			10709 => std_logic_vector(to_unsigned( 151,8)),
			10710 => std_logic_vector(to_unsigned( 124,8)),
			10711 => std_logic_vector(to_unsigned( 246,8)),
			10712 => std_logic_vector(to_unsigned( 246,8)),
			10713 => std_logic_vector(to_unsigned( 180,8)),
			10714 => std_logic_vector(to_unsigned( 148,8)),
			10715 => std_logic_vector(to_unsigned( 134,8)),
			10716 => std_logic_vector(to_unsigned( 79,8)),
			10717 => std_logic_vector(to_unsigned( 144,8)),
			10718 => std_logic_vector(to_unsigned( 7,8)),
			10719 => std_logic_vector(to_unsigned( 229,8)),
			10720 => std_logic_vector(to_unsigned( 197,8)),
			10721 => std_logic_vector(to_unsigned( 104,8)),
			10722 => std_logic_vector(to_unsigned( 130,8)),
			10723 => std_logic_vector(to_unsigned( 104,8)),
			10724 => std_logic_vector(to_unsigned( 65,8)),
			10725 => std_logic_vector(to_unsigned( 98,8)),
			10726 => std_logic_vector(to_unsigned( 236,8)),
			10727 => std_logic_vector(to_unsigned( 139,8)),
			10728 => std_logic_vector(to_unsigned( 74,8)),
			10729 => std_logic_vector(to_unsigned( 41,8)),
			10730 => std_logic_vector(to_unsigned( 146,8)),
			10731 => std_logic_vector(to_unsigned( 35,8)),
			10732 => std_logic_vector(to_unsigned( 89,8)),
			10733 => std_logic_vector(to_unsigned( 137,8)),
			10734 => std_logic_vector(to_unsigned( 223,8)),
			10735 => std_logic_vector(to_unsigned( 63,8)),
			10736 => std_logic_vector(to_unsigned( 193,8)),
			10737 => std_logic_vector(to_unsigned( 160,8)),
			10738 => std_logic_vector(to_unsigned( 18,8)),
			10739 => std_logic_vector(to_unsigned( 120,8)),
			10740 => std_logic_vector(to_unsigned( 250,8)),
			10741 => std_logic_vector(to_unsigned( 146,8)),
			10742 => std_logic_vector(to_unsigned( 238,8)),
			10743 => std_logic_vector(to_unsigned( 227,8)),
			10744 => std_logic_vector(to_unsigned( 128,8)),
			10745 => std_logic_vector(to_unsigned( 250,8)),
			10746 => std_logic_vector(to_unsigned( 234,8)),
			10747 => std_logic_vector(to_unsigned( 157,8)),
			10748 => std_logic_vector(to_unsigned( 122,8)),
			10749 => std_logic_vector(to_unsigned( 39,8)),
			10750 => std_logic_vector(to_unsigned( 111,8)),
			10751 => std_logic_vector(to_unsigned( 137,8)),
			10752 => std_logic_vector(to_unsigned( 125,8)),
			10753 => std_logic_vector(to_unsigned( 41,8)),
			10754 => std_logic_vector(to_unsigned( 231,8)),
			10755 => std_logic_vector(to_unsigned( 106,8)),
			10756 => std_logic_vector(to_unsigned( 96,8)),
			10757 => std_logic_vector(to_unsigned( 241,8)),
			10758 => std_logic_vector(to_unsigned( 47,8)),
			10759 => std_logic_vector(to_unsigned( 246,8)),
			10760 => std_logic_vector(to_unsigned( 130,8)),
			10761 => std_logic_vector(to_unsigned( 89,8)),
			10762 => std_logic_vector(to_unsigned( 44,8)),
			10763 => std_logic_vector(to_unsigned( 118,8)),
			10764 => std_logic_vector(to_unsigned( 69,8)),
			10765 => std_logic_vector(to_unsigned( 25,8)),
			10766 => std_logic_vector(to_unsigned( 54,8)),
			10767 => std_logic_vector(to_unsigned( 171,8)),
			10768 => std_logic_vector(to_unsigned( 61,8)),
			10769 => std_logic_vector(to_unsigned( 80,8)),
			10770 => std_logic_vector(to_unsigned( 49,8)),
			10771 => std_logic_vector(to_unsigned( 105,8)),
			10772 => std_logic_vector(to_unsigned( 171,8)),
			10773 => std_logic_vector(to_unsigned( 116,8)),
			10774 => std_logic_vector(to_unsigned( 83,8)),
			10775 => std_logic_vector(to_unsigned( 152,8)),
			10776 => std_logic_vector(to_unsigned( 62,8)),
			10777 => std_logic_vector(to_unsigned( 90,8)),
			10778 => std_logic_vector(to_unsigned( 44,8)),
			10779 => std_logic_vector(to_unsigned( 60,8)),
			10780 => std_logic_vector(to_unsigned( 95,8)),
			10781 => std_logic_vector(to_unsigned( 32,8)),
			10782 => std_logic_vector(to_unsigned( 108,8)),
			10783 => std_logic_vector(to_unsigned( 6,8)),
			10784 => std_logic_vector(to_unsigned( 223,8)),
			10785 => std_logic_vector(to_unsigned( 83,8)),
			10786 => std_logic_vector(to_unsigned( 84,8)),
			10787 => std_logic_vector(to_unsigned( 18,8)),
			10788 => std_logic_vector(to_unsigned( 89,8)),
			10789 => std_logic_vector(to_unsigned( 80,8)),
			10790 => std_logic_vector(to_unsigned( 10,8)),
			10791 => std_logic_vector(to_unsigned( 151,8)),
			10792 => std_logic_vector(to_unsigned( 245,8)),
			10793 => std_logic_vector(to_unsigned( 225,8)),
			10794 => std_logic_vector(to_unsigned( 29,8)),
			10795 => std_logic_vector(to_unsigned( 230,8)),
			10796 => std_logic_vector(to_unsigned( 189,8)),
			10797 => std_logic_vector(to_unsigned( 46,8)),
			10798 => std_logic_vector(to_unsigned( 15,8)),
			10799 => std_logic_vector(to_unsigned( 20,8)),
			10800 => std_logic_vector(to_unsigned( 250,8)),
			10801 => std_logic_vector(to_unsigned( 97,8)),
			10802 => std_logic_vector(to_unsigned( 87,8)),
			10803 => std_logic_vector(to_unsigned( 188,8)),
			10804 => std_logic_vector(to_unsigned( 189,8)),
			10805 => std_logic_vector(to_unsigned( 30,8)),
			10806 => std_logic_vector(to_unsigned( 103,8)),
			10807 => std_logic_vector(to_unsigned( 58,8)),
			10808 => std_logic_vector(to_unsigned( 232,8)),
			10809 => std_logic_vector(to_unsigned( 218,8)),
			10810 => std_logic_vector(to_unsigned( 188,8)),
			10811 => std_logic_vector(to_unsigned( 190,8)),
			10812 => std_logic_vector(to_unsigned( 96,8)),
			10813 => std_logic_vector(to_unsigned( 224,8)),
			10814 => std_logic_vector(to_unsigned( 196,8)),
			10815 => std_logic_vector(to_unsigned( 177,8)),
			10816 => std_logic_vector(to_unsigned( 60,8)),
			10817 => std_logic_vector(to_unsigned( 158,8)),
			10818 => std_logic_vector(to_unsigned( 136,8)),
			10819 => std_logic_vector(to_unsigned( 183,8)),
			10820 => std_logic_vector(to_unsigned( 21,8)),
			10821 => std_logic_vector(to_unsigned( 153,8)),
			10822 => std_logic_vector(to_unsigned( 97,8)),
			10823 => std_logic_vector(to_unsigned( 202,8)),
			10824 => std_logic_vector(to_unsigned( 50,8)),
			10825 => std_logic_vector(to_unsigned( 180,8)),
			10826 => std_logic_vector(to_unsigned( 94,8)),
			10827 => std_logic_vector(to_unsigned( 247,8)),
			10828 => std_logic_vector(to_unsigned( 236,8)),
			10829 => std_logic_vector(to_unsigned( 34,8)),
			10830 => std_logic_vector(to_unsigned( 150,8)),
			10831 => std_logic_vector(to_unsigned( 178,8)),
			10832 => std_logic_vector(to_unsigned( 122,8)),
			10833 => std_logic_vector(to_unsigned( 70,8)),
			10834 => std_logic_vector(to_unsigned( 194,8)),
			10835 => std_logic_vector(to_unsigned( 43,8)),
			10836 => std_logic_vector(to_unsigned( 18,8)),
			10837 => std_logic_vector(to_unsigned( 226,8)),
			10838 => std_logic_vector(to_unsigned( 50,8)),
			10839 => std_logic_vector(to_unsigned( 141,8)),
			10840 => std_logic_vector(to_unsigned( 189,8)),
			10841 => std_logic_vector(to_unsigned( 104,8)),
			10842 => std_logic_vector(to_unsigned( 192,8)),
			10843 => std_logic_vector(to_unsigned( 67,8)),
			10844 => std_logic_vector(to_unsigned( 93,8)),
			10845 => std_logic_vector(to_unsigned( 159,8)),
			10846 => std_logic_vector(to_unsigned( 46,8)),
			10847 => std_logic_vector(to_unsigned( 45,8)),
			10848 => std_logic_vector(to_unsigned( 20,8)),
			10849 => std_logic_vector(to_unsigned( 22,8)),
			10850 => std_logic_vector(to_unsigned( 40,8)),
			10851 => std_logic_vector(to_unsigned( 6,8)),
			10852 => std_logic_vector(to_unsigned( 237,8)),
			10853 => std_logic_vector(to_unsigned( 70,8)),
			10854 => std_logic_vector(to_unsigned( 247,8)),
			10855 => std_logic_vector(to_unsigned( 92,8)),
			10856 => std_logic_vector(to_unsigned( 104,8)),
			10857 => std_logic_vector(to_unsigned( 99,8)),
			10858 => std_logic_vector(to_unsigned( 98,8)),
			10859 => std_logic_vector(to_unsigned( 236,8)),
			10860 => std_logic_vector(to_unsigned( 255,8)),
			10861 => std_logic_vector(to_unsigned( 53,8)),
			10862 => std_logic_vector(to_unsigned( 83,8)),
			10863 => std_logic_vector(to_unsigned( 196,8)),
			10864 => std_logic_vector(to_unsigned( 112,8)),
			10865 => std_logic_vector(to_unsigned( 133,8)),
			10866 => std_logic_vector(to_unsigned( 94,8)),
			10867 => std_logic_vector(to_unsigned( 199,8)),
			10868 => std_logic_vector(to_unsigned( 105,8)),
			10869 => std_logic_vector(to_unsigned( 56,8)),
			10870 => std_logic_vector(to_unsigned( 224,8)),
			10871 => std_logic_vector(to_unsigned( 73,8)),
			10872 => std_logic_vector(to_unsigned( 237,8)),
			10873 => std_logic_vector(to_unsigned( 179,8)),
			10874 => std_logic_vector(to_unsigned( 228,8)),
			10875 => std_logic_vector(to_unsigned( 85,8)),
			10876 => std_logic_vector(to_unsigned( 230,8)),
			10877 => std_logic_vector(to_unsigned( 225,8)),
			10878 => std_logic_vector(to_unsigned( 219,8)),
			10879 => std_logic_vector(to_unsigned( 85,8)),
			10880 => std_logic_vector(to_unsigned( 167,8)),
			10881 => std_logic_vector(to_unsigned( 192,8)),
			10882 => std_logic_vector(to_unsigned( 41,8)),
			10883 => std_logic_vector(to_unsigned( 194,8)),
			10884 => std_logic_vector(to_unsigned( 248,8)),
			10885 => std_logic_vector(to_unsigned( 167,8)),
			10886 => std_logic_vector(to_unsigned( 176,8)),
			10887 => std_logic_vector(to_unsigned( 37,8)),
			10888 => std_logic_vector(to_unsigned( 3,8)),
			10889 => std_logic_vector(to_unsigned( 182,8)),
			10890 => std_logic_vector(to_unsigned( 84,8)),
			10891 => std_logic_vector(to_unsigned( 31,8)),
			10892 => std_logic_vector(to_unsigned( 154,8)),
			10893 => std_logic_vector(to_unsigned( 81,8)),
			10894 => std_logic_vector(to_unsigned( 221,8)),
			10895 => std_logic_vector(to_unsigned( 60,8)),
			10896 => std_logic_vector(to_unsigned( 59,8)),
			10897 => std_logic_vector(to_unsigned( 132,8)),
			10898 => std_logic_vector(to_unsigned( 241,8)),
			10899 => std_logic_vector(to_unsigned( 235,8)),
			10900 => std_logic_vector(to_unsigned( 146,8)),
			10901 => std_logic_vector(to_unsigned( 125,8)),
			10902 => std_logic_vector(to_unsigned( 206,8)),
			10903 => std_logic_vector(to_unsigned( 68,8)),
			10904 => std_logic_vector(to_unsigned( 26,8)),
			10905 => std_logic_vector(to_unsigned( 58,8)),
			10906 => std_logic_vector(to_unsigned( 131,8)),
			10907 => std_logic_vector(to_unsigned( 231,8)),
			10908 => std_logic_vector(to_unsigned( 172,8)),
			10909 => std_logic_vector(to_unsigned( 248,8)),
			10910 => std_logic_vector(to_unsigned( 214,8)),
			10911 => std_logic_vector(to_unsigned( 57,8)),
			10912 => std_logic_vector(to_unsigned( 43,8)),
			10913 => std_logic_vector(to_unsigned( 79,8)),
			10914 => std_logic_vector(to_unsigned( 250,8)),
			10915 => std_logic_vector(to_unsigned( 233,8)),
			10916 => std_logic_vector(to_unsigned( 199,8)),
			10917 => std_logic_vector(to_unsigned( 154,8)),
			10918 => std_logic_vector(to_unsigned( 40,8)),
			10919 => std_logic_vector(to_unsigned( 245,8)),
			10920 => std_logic_vector(to_unsigned( 168,8)),
			10921 => std_logic_vector(to_unsigned( 36,8)),
			10922 => std_logic_vector(to_unsigned( 72,8)),
			10923 => std_logic_vector(to_unsigned( 67,8)),
			10924 => std_logic_vector(to_unsigned( 11,8)),
			10925 => std_logic_vector(to_unsigned( 100,8)),
			10926 => std_logic_vector(to_unsigned( 142,8)),
			10927 => std_logic_vector(to_unsigned( 186,8)),
			10928 => std_logic_vector(to_unsigned( 89,8)),
			10929 => std_logic_vector(to_unsigned( 194,8)),
			10930 => std_logic_vector(to_unsigned( 78,8)),
			10931 => std_logic_vector(to_unsigned( 58,8)),
			10932 => std_logic_vector(to_unsigned( 221,8)),
			10933 => std_logic_vector(to_unsigned( 30,8)),
			10934 => std_logic_vector(to_unsigned( 236,8)),
			10935 => std_logic_vector(to_unsigned( 114,8)),
			10936 => std_logic_vector(to_unsigned( 167,8)),
			10937 => std_logic_vector(to_unsigned( 74,8)),
			10938 => std_logic_vector(to_unsigned( 50,8)),
			10939 => std_logic_vector(to_unsigned( 159,8)),
			10940 => std_logic_vector(to_unsigned( 160,8)),
			10941 => std_logic_vector(to_unsigned( 107,8)),
			10942 => std_logic_vector(to_unsigned( 79,8)),
			10943 => std_logic_vector(to_unsigned( 2,8)),
			10944 => std_logic_vector(to_unsigned( 14,8)),
			10945 => std_logic_vector(to_unsigned( 3,8)),
			10946 => std_logic_vector(to_unsigned( 114,8)),
			10947 => std_logic_vector(to_unsigned( 67,8)),
			10948 => std_logic_vector(to_unsigned( 168,8)),
			10949 => std_logic_vector(to_unsigned( 22,8)),
			10950 => std_logic_vector(to_unsigned( 218,8)),
			10951 => std_logic_vector(to_unsigned( 29,8)),
			10952 => std_logic_vector(to_unsigned( 41,8)),
			10953 => std_logic_vector(to_unsigned( 25,8)),
			10954 => std_logic_vector(to_unsigned( 208,8)),
			10955 => std_logic_vector(to_unsigned( 199,8)),
			10956 => std_logic_vector(to_unsigned( 112,8)),
			10957 => std_logic_vector(to_unsigned( 247,8)),
			10958 => std_logic_vector(to_unsigned( 65,8)),
			10959 => std_logic_vector(to_unsigned( 144,8)),
			10960 => std_logic_vector(to_unsigned( 88,8)),
			10961 => std_logic_vector(to_unsigned( 50,8)),
			10962 => std_logic_vector(to_unsigned( 141,8)),
			10963 => std_logic_vector(to_unsigned( 29,8)),
			10964 => std_logic_vector(to_unsigned( 250,8)),
			10965 => std_logic_vector(to_unsigned( 144,8)),
			10966 => std_logic_vector(to_unsigned( 44,8)),
			10967 => std_logic_vector(to_unsigned( 180,8)),
			10968 => std_logic_vector(to_unsigned( 234,8)),
			10969 => std_logic_vector(to_unsigned( 201,8)),
			10970 => std_logic_vector(to_unsigned( 97,8)),
			10971 => std_logic_vector(to_unsigned( 136,8)),
			10972 => std_logic_vector(to_unsigned( 0,8)),
			10973 => std_logic_vector(to_unsigned( 167,8)),
			10974 => std_logic_vector(to_unsigned( 245,8)),
			10975 => std_logic_vector(to_unsigned( 5,8)),
			10976 => std_logic_vector(to_unsigned( 142,8)),
			10977 => std_logic_vector(to_unsigned( 153,8)),
			10978 => std_logic_vector(to_unsigned( 34,8)),
			10979 => std_logic_vector(to_unsigned( 35,8)),
			10980 => std_logic_vector(to_unsigned( 146,8)),
			10981 => std_logic_vector(to_unsigned( 138,8)),
			10982 => std_logic_vector(to_unsigned( 113,8)),
			10983 => std_logic_vector(to_unsigned( 88,8)),
			10984 => std_logic_vector(to_unsigned( 230,8)),
			10985 => std_logic_vector(to_unsigned( 237,8)),
			10986 => std_logic_vector(to_unsigned( 206,8)),
			10987 => std_logic_vector(to_unsigned( 165,8)),
			10988 => std_logic_vector(to_unsigned( 245,8)),
			10989 => std_logic_vector(to_unsigned( 50,8)),
			10990 => std_logic_vector(to_unsigned( 156,8)),
			10991 => std_logic_vector(to_unsigned( 189,8)),
			10992 => std_logic_vector(to_unsigned( 235,8)),
			10993 => std_logic_vector(to_unsigned( 52,8)),
			10994 => std_logic_vector(to_unsigned( 64,8)),
			10995 => std_logic_vector(to_unsigned( 21,8)),
			10996 => std_logic_vector(to_unsigned( 28,8)),
			10997 => std_logic_vector(to_unsigned( 156,8)),
			10998 => std_logic_vector(to_unsigned( 212,8)),
			10999 => std_logic_vector(to_unsigned( 130,8)),
			11000 => std_logic_vector(to_unsigned( 118,8)),
			11001 => std_logic_vector(to_unsigned( 129,8)),
			11002 => std_logic_vector(to_unsigned( 142,8)),
			11003 => std_logic_vector(to_unsigned( 91,8)),
			11004 => std_logic_vector(to_unsigned( 18,8)),
			11005 => std_logic_vector(to_unsigned( 28,8)),
			11006 => std_logic_vector(to_unsigned( 118,8)),
			11007 => std_logic_vector(to_unsigned( 208,8)),
			11008 => std_logic_vector(to_unsigned( 146,8)),
			11009 => std_logic_vector(to_unsigned( 160,8)),
			11010 => std_logic_vector(to_unsigned( 220,8)),
			11011 => std_logic_vector(to_unsigned( 167,8)),
			11012 => std_logic_vector(to_unsigned( 142,8)),
			11013 => std_logic_vector(to_unsigned( 141,8)),
			11014 => std_logic_vector(to_unsigned( 223,8)),
			11015 => std_logic_vector(to_unsigned( 212,8)),
			11016 => std_logic_vector(to_unsigned( 129,8)),
			11017 => std_logic_vector(to_unsigned( 3,8)),
			11018 => std_logic_vector(to_unsigned( 222,8)),
			11019 => std_logic_vector(to_unsigned( 227,8)),
			11020 => std_logic_vector(to_unsigned( 245,8)),
			11021 => std_logic_vector(to_unsigned( 63,8)),
			11022 => std_logic_vector(to_unsigned( 13,8)),
			11023 => std_logic_vector(to_unsigned( 64,8)),
			11024 => std_logic_vector(to_unsigned( 249,8)),
			11025 => std_logic_vector(to_unsigned( 253,8)),
			11026 => std_logic_vector(to_unsigned( 118,8)),
			11027 => std_logic_vector(to_unsigned( 8,8)),
			11028 => std_logic_vector(to_unsigned( 20,8)),
			11029 => std_logic_vector(to_unsigned( 26,8)),
			11030 => std_logic_vector(to_unsigned( 76,8)),
			11031 => std_logic_vector(to_unsigned( 248,8)),
			11032 => std_logic_vector(to_unsigned( 119,8)),
			11033 => std_logic_vector(to_unsigned( 75,8)),
			11034 => std_logic_vector(to_unsigned( 210,8)),
			11035 => std_logic_vector(to_unsigned( 201,8)),
			11036 => std_logic_vector(to_unsigned( 214,8)),
			11037 => std_logic_vector(to_unsigned( 230,8)),
			11038 => std_logic_vector(to_unsigned( 31,8)),
			11039 => std_logic_vector(to_unsigned( 103,8)),
			11040 => std_logic_vector(to_unsigned( 187,8)),
			11041 => std_logic_vector(to_unsigned( 225,8)),
			11042 => std_logic_vector(to_unsigned( 5,8)),
			11043 => std_logic_vector(to_unsigned( 19,8)),
			11044 => std_logic_vector(to_unsigned( 95,8)),
			11045 => std_logic_vector(to_unsigned( 18,8)),
			11046 => std_logic_vector(to_unsigned( 208,8)),
			11047 => std_logic_vector(to_unsigned( 118,8)),
			11048 => std_logic_vector(to_unsigned( 171,8)),
			11049 => std_logic_vector(to_unsigned( 69,8)),
			11050 => std_logic_vector(to_unsigned( 45,8)),
			11051 => std_logic_vector(to_unsigned( 143,8)),
			11052 => std_logic_vector(to_unsigned( 141,8)),
			11053 => std_logic_vector(to_unsigned( 53,8)),
			11054 => std_logic_vector(to_unsigned( 75,8)),
			11055 => std_logic_vector(to_unsigned( 224,8)),
			11056 => std_logic_vector(to_unsigned( 178,8)),
			11057 => std_logic_vector(to_unsigned( 36,8)),
			11058 => std_logic_vector(to_unsigned( 54,8)),
			11059 => std_logic_vector(to_unsigned( 8,8)),
			11060 => std_logic_vector(to_unsigned( 13,8)),
			11061 => std_logic_vector(to_unsigned( 248,8)),
			11062 => std_logic_vector(to_unsigned( 196,8)),
			11063 => std_logic_vector(to_unsigned( 14,8)),
			11064 => std_logic_vector(to_unsigned( 225,8)),
			11065 => std_logic_vector(to_unsigned( 24,8)),
			11066 => std_logic_vector(to_unsigned( 229,8)),
			11067 => std_logic_vector(to_unsigned( 53,8)),
			11068 => std_logic_vector(to_unsigned( 32,8)),
			11069 => std_logic_vector(to_unsigned( 190,8)),
			11070 => std_logic_vector(to_unsigned( 33,8)),
			11071 => std_logic_vector(to_unsigned( 71,8)),
			11072 => std_logic_vector(to_unsigned( 204,8)),
			11073 => std_logic_vector(to_unsigned( 221,8)),
			11074 => std_logic_vector(to_unsigned( 239,8)),
			11075 => std_logic_vector(to_unsigned( 192,8)),
			11076 => std_logic_vector(to_unsigned( 148,8)),
			11077 => std_logic_vector(to_unsigned( 195,8)),
			11078 => std_logic_vector(to_unsigned( 199,8)),
			11079 => std_logic_vector(to_unsigned( 7,8)),
			11080 => std_logic_vector(to_unsigned( 3,8)),
			11081 => std_logic_vector(to_unsigned( 82,8)),
			11082 => std_logic_vector(to_unsigned( 199,8)),
			11083 => std_logic_vector(to_unsigned( 196,8)),
			11084 => std_logic_vector(to_unsigned( 147,8)),
			11085 => std_logic_vector(to_unsigned( 92,8)),
			11086 => std_logic_vector(to_unsigned( 140,8)),
			11087 => std_logic_vector(to_unsigned( 63,8)),
			11088 => std_logic_vector(to_unsigned( 8,8)),
			11089 => std_logic_vector(to_unsigned( 75,8)),
			11090 => std_logic_vector(to_unsigned( 119,8)),
			11091 => std_logic_vector(to_unsigned( 136,8)),
			11092 => std_logic_vector(to_unsigned( 71,8)),
			11093 => std_logic_vector(to_unsigned( 8,8)),
			11094 => std_logic_vector(to_unsigned( 203,8)),
			11095 => std_logic_vector(to_unsigned( 236,8)),
			11096 => std_logic_vector(to_unsigned( 163,8)),
			11097 => std_logic_vector(to_unsigned( 184,8)),
			11098 => std_logic_vector(to_unsigned( 145,8)),
			11099 => std_logic_vector(to_unsigned( 88,8)),
			11100 => std_logic_vector(to_unsigned( 47,8)),
			11101 => std_logic_vector(to_unsigned( 26,8)),
			11102 => std_logic_vector(to_unsigned( 61,8)),
			11103 => std_logic_vector(to_unsigned( 245,8)),
			11104 => std_logic_vector(to_unsigned( 79,8)),
			11105 => std_logic_vector(to_unsigned( 222,8)),
			11106 => std_logic_vector(to_unsigned( 76,8)),
			11107 => std_logic_vector(to_unsigned( 112,8)),
			11108 => std_logic_vector(to_unsigned( 143,8)),
			11109 => std_logic_vector(to_unsigned( 184,8)),
			11110 => std_logic_vector(to_unsigned( 51,8)),
			11111 => std_logic_vector(to_unsigned( 107,8)),
			11112 => std_logic_vector(to_unsigned( 250,8)),
			11113 => std_logic_vector(to_unsigned( 101,8)),
			11114 => std_logic_vector(to_unsigned( 40,8)),
			11115 => std_logic_vector(to_unsigned( 181,8)),
			11116 => std_logic_vector(to_unsigned( 121,8)),
			11117 => std_logic_vector(to_unsigned( 51,8)),
			11118 => std_logic_vector(to_unsigned( 6,8)),
			11119 => std_logic_vector(to_unsigned( 219,8)),
			11120 => std_logic_vector(to_unsigned( 154,8)),
			11121 => std_logic_vector(to_unsigned( 28,8)),
			11122 => std_logic_vector(to_unsigned( 65,8)),
			11123 => std_logic_vector(to_unsigned( 138,8)),
			11124 => std_logic_vector(to_unsigned( 233,8)),
			11125 => std_logic_vector(to_unsigned( 137,8)),
			11126 => std_logic_vector(to_unsigned( 212,8)),
			11127 => std_logic_vector(to_unsigned( 196,8)),
			11128 => std_logic_vector(to_unsigned( 245,8)),
			11129 => std_logic_vector(to_unsigned( 93,8)),
			11130 => std_logic_vector(to_unsigned( 135,8)),
			11131 => std_logic_vector(to_unsigned( 3,8)),
			11132 => std_logic_vector(to_unsigned( 47,8)),
			11133 => std_logic_vector(to_unsigned( 45,8)),
			11134 => std_logic_vector(to_unsigned( 212,8)),
			11135 => std_logic_vector(to_unsigned( 51,8)),
			11136 => std_logic_vector(to_unsigned( 245,8)),
			11137 => std_logic_vector(to_unsigned( 82,8)),
			11138 => std_logic_vector(to_unsigned( 220,8)),
			11139 => std_logic_vector(to_unsigned( 239,8)),
			11140 => std_logic_vector(to_unsigned( 132,8)),
			11141 => std_logic_vector(to_unsigned( 80,8)),
			11142 => std_logic_vector(to_unsigned( 126,8)),
			11143 => std_logic_vector(to_unsigned( 208,8)),
			11144 => std_logic_vector(to_unsigned( 65,8)),
			11145 => std_logic_vector(to_unsigned( 122,8)),
			11146 => std_logic_vector(to_unsigned( 235,8)),
			11147 => std_logic_vector(to_unsigned( 70,8)),
			11148 => std_logic_vector(to_unsigned( 134,8)),
			11149 => std_logic_vector(to_unsigned( 23,8)),
			11150 => std_logic_vector(to_unsigned( 115,8)),
			11151 => std_logic_vector(to_unsigned( 0,8)),
			11152 => std_logic_vector(to_unsigned( 91,8)),
			11153 => std_logic_vector(to_unsigned( 56,8)),
			11154 => std_logic_vector(to_unsigned( 239,8)),
			11155 => std_logic_vector(to_unsigned( 95,8)),
			11156 => std_logic_vector(to_unsigned( 129,8)),
			11157 => std_logic_vector(to_unsigned( 89,8)),
			11158 => std_logic_vector(to_unsigned( 51,8)),
			11159 => std_logic_vector(to_unsigned( 226,8)),
			11160 => std_logic_vector(to_unsigned( 152,8)),
			11161 => std_logic_vector(to_unsigned( 25,8)),
			11162 => std_logic_vector(to_unsigned( 164,8)),
			11163 => std_logic_vector(to_unsigned( 190,8)),
			11164 => std_logic_vector(to_unsigned( 242,8)),
			11165 => std_logic_vector(to_unsigned( 7,8)),
			11166 => std_logic_vector(to_unsigned( 29,8)),
			11167 => std_logic_vector(to_unsigned( 172,8)),
			11168 => std_logic_vector(to_unsigned( 183,8)),
			11169 => std_logic_vector(to_unsigned( 152,8)),
			11170 => std_logic_vector(to_unsigned( 30,8)),
			11171 => std_logic_vector(to_unsigned( 136,8)),
			11172 => std_logic_vector(to_unsigned( 91,8)),
			11173 => std_logic_vector(to_unsigned( 164,8)),
			11174 => std_logic_vector(to_unsigned( 106,8)),
			11175 => std_logic_vector(to_unsigned( 187,8)),
			11176 => std_logic_vector(to_unsigned( 70,8)),
			11177 => std_logic_vector(to_unsigned( 125,8)),
			11178 => std_logic_vector(to_unsigned( 165,8)),
			11179 => std_logic_vector(to_unsigned( 225,8)),
			11180 => std_logic_vector(to_unsigned( 191,8)),
			11181 => std_logic_vector(to_unsigned( 50,8)),
			11182 => std_logic_vector(to_unsigned( 82,8)),
			11183 => std_logic_vector(to_unsigned( 150,8)),
			11184 => std_logic_vector(to_unsigned( 6,8)),
			11185 => std_logic_vector(to_unsigned( 119,8)),
			11186 => std_logic_vector(to_unsigned( 227,8)),
			11187 => std_logic_vector(to_unsigned( 44,8)),
			11188 => std_logic_vector(to_unsigned( 250,8)),
			11189 => std_logic_vector(to_unsigned( 96,8)),
			11190 => std_logic_vector(to_unsigned( 98,8)),
			11191 => std_logic_vector(to_unsigned( 60,8)),
			11192 => std_logic_vector(to_unsigned( 79,8)),
			11193 => std_logic_vector(to_unsigned( 213,8)),
			11194 => std_logic_vector(to_unsigned( 126,8)),
			11195 => std_logic_vector(to_unsigned( 2,8)),
			11196 => std_logic_vector(to_unsigned( 59,8)),
			11197 => std_logic_vector(to_unsigned( 26,8)),
			11198 => std_logic_vector(to_unsigned( 222,8)),
			11199 => std_logic_vector(to_unsigned( 99,8)),
			11200 => std_logic_vector(to_unsigned( 31,8)),
			11201 => std_logic_vector(to_unsigned( 178,8)),
			11202 => std_logic_vector(to_unsigned( 229,8)),
			11203 => std_logic_vector(to_unsigned( 76,8)),
			11204 => std_logic_vector(to_unsigned( 137,8)),
			11205 => std_logic_vector(to_unsigned( 29,8)),
			11206 => std_logic_vector(to_unsigned( 4,8)),
			11207 => std_logic_vector(to_unsigned( 129,8)),
			11208 => std_logic_vector(to_unsigned( 52,8)),
			11209 => std_logic_vector(to_unsigned( 11,8)),
			11210 => std_logic_vector(to_unsigned( 191,8)),
			11211 => std_logic_vector(to_unsigned( 56,8)),
			11212 => std_logic_vector(to_unsigned( 119,8)),
			11213 => std_logic_vector(to_unsigned( 232,8)),
			11214 => std_logic_vector(to_unsigned( 28,8)),
			11215 => std_logic_vector(to_unsigned( 136,8)),
			11216 => std_logic_vector(to_unsigned( 245,8)),
			11217 => std_logic_vector(to_unsigned( 28,8)),
			11218 => std_logic_vector(to_unsigned( 119,8)),
			11219 => std_logic_vector(to_unsigned( 76,8)),
			11220 => std_logic_vector(to_unsigned( 62,8)),
			11221 => std_logic_vector(to_unsigned( 145,8)),
			11222 => std_logic_vector(to_unsigned( 231,8)),
			11223 => std_logic_vector(to_unsigned( 29,8)),
			11224 => std_logic_vector(to_unsigned( 86,8)),
			11225 => std_logic_vector(to_unsigned( 235,8)),
			11226 => std_logic_vector(to_unsigned( 204,8)),
			11227 => std_logic_vector(to_unsigned( 47,8)),
			11228 => std_logic_vector(to_unsigned( 227,8)),
			11229 => std_logic_vector(to_unsigned( 93,8)),
			11230 => std_logic_vector(to_unsigned( 102,8)),
			11231 => std_logic_vector(to_unsigned( 82,8)),
			11232 => std_logic_vector(to_unsigned( 116,8)),
			11233 => std_logic_vector(to_unsigned( 13,8)),
			11234 => std_logic_vector(to_unsigned( 88,8)),
			11235 => std_logic_vector(to_unsigned( 213,8)),
			11236 => std_logic_vector(to_unsigned( 247,8)),
			11237 => std_logic_vector(to_unsigned( 37,8)),
			11238 => std_logic_vector(to_unsigned( 198,8)),
			11239 => std_logic_vector(to_unsigned( 122,8)),
			11240 => std_logic_vector(to_unsigned( 151,8)),
			11241 => std_logic_vector(to_unsigned( 198,8)),
			11242 => std_logic_vector(to_unsigned( 218,8)),
			11243 => std_logic_vector(to_unsigned( 35,8)),
			11244 => std_logic_vector(to_unsigned( 83,8)),
			11245 => std_logic_vector(to_unsigned( 12,8)),
			11246 => std_logic_vector(to_unsigned( 20,8)),
			11247 => std_logic_vector(to_unsigned( 234,8)),
			11248 => std_logic_vector(to_unsigned( 98,8)),
			11249 => std_logic_vector(to_unsigned( 127,8)),
			11250 => std_logic_vector(to_unsigned( 62,8)),
			11251 => std_logic_vector(to_unsigned( 127,8)),
			11252 => std_logic_vector(to_unsigned( 100,8)),
			11253 => std_logic_vector(to_unsigned( 232,8)),
			11254 => std_logic_vector(to_unsigned( 25,8)),
			11255 => std_logic_vector(to_unsigned( 239,8)),
			11256 => std_logic_vector(to_unsigned( 121,8)),
			11257 => std_logic_vector(to_unsigned( 51,8)),
			11258 => std_logic_vector(to_unsigned( 215,8)),
			11259 => std_logic_vector(to_unsigned( 222,8)),
			11260 => std_logic_vector(to_unsigned( 3,8)),
			11261 => std_logic_vector(to_unsigned( 30,8)),
			11262 => std_logic_vector(to_unsigned( 99,8)),
			11263 => std_logic_vector(to_unsigned( 214,8)),
			11264 => std_logic_vector(to_unsigned( 123,8)),
			11265 => std_logic_vector(to_unsigned( 112,8)),
			11266 => std_logic_vector(to_unsigned( 159,8)),
			11267 => std_logic_vector(to_unsigned( 116,8)),
			11268 => std_logic_vector(to_unsigned( 197,8)),
			11269 => std_logic_vector(to_unsigned( 74,8)),
			11270 => std_logic_vector(to_unsigned( 15,8)),
			11271 => std_logic_vector(to_unsigned( 31,8)),
			11272 => std_logic_vector(to_unsigned( 189,8)),
			11273 => std_logic_vector(to_unsigned( 7,8)),
			11274 => std_logic_vector(to_unsigned( 254,8)),
			11275 => std_logic_vector(to_unsigned( 195,8)),
			11276 => std_logic_vector(to_unsigned( 108,8)),
			11277 => std_logic_vector(to_unsigned( 35,8)),
			11278 => std_logic_vector(to_unsigned( 246,8)),
			11279 => std_logic_vector(to_unsigned( 124,8)),
			11280 => std_logic_vector(to_unsigned( 251,8)),
			11281 => std_logic_vector(to_unsigned( 82,8)),
			11282 => std_logic_vector(to_unsigned( 61,8)),
			11283 => std_logic_vector(to_unsigned( 121,8)),
			11284 => std_logic_vector(to_unsigned( 99,8)),
			11285 => std_logic_vector(to_unsigned( 106,8)),
			11286 => std_logic_vector(to_unsigned( 143,8)),
			11287 => std_logic_vector(to_unsigned( 235,8)),
			11288 => std_logic_vector(to_unsigned( 96,8)),
			11289 => std_logic_vector(to_unsigned( 192,8)),
			11290 => std_logic_vector(to_unsigned( 253,8)),
			11291 => std_logic_vector(to_unsigned( 138,8)),
			11292 => std_logic_vector(to_unsigned( 41,8)),
			11293 => std_logic_vector(to_unsigned( 198,8)),
			11294 => std_logic_vector(to_unsigned( 217,8)),
			11295 => std_logic_vector(to_unsigned( 46,8)),
			11296 => std_logic_vector(to_unsigned( 117,8)),
			11297 => std_logic_vector(to_unsigned( 206,8)),
			11298 => std_logic_vector(to_unsigned( 102,8)),
			11299 => std_logic_vector(to_unsigned( 67,8)),
			11300 => std_logic_vector(to_unsigned( 199,8)),
			11301 => std_logic_vector(to_unsigned( 142,8)),
			11302 => std_logic_vector(to_unsigned( 240,8)),
			11303 => std_logic_vector(to_unsigned( 20,8)),
			11304 => std_logic_vector(to_unsigned( 129,8)),
			11305 => std_logic_vector(to_unsigned( 50,8)),
			11306 => std_logic_vector(to_unsigned( 231,8)),
			11307 => std_logic_vector(to_unsigned( 12,8)),
			11308 => std_logic_vector(to_unsigned( 174,8)),
			11309 => std_logic_vector(to_unsigned( 63,8)),
			11310 => std_logic_vector(to_unsigned( 210,8)),
			11311 => std_logic_vector(to_unsigned( 162,8)),
			11312 => std_logic_vector(to_unsigned( 10,8)),
			11313 => std_logic_vector(to_unsigned( 25,8)),
			11314 => std_logic_vector(to_unsigned( 85,8)),
			11315 => std_logic_vector(to_unsigned( 103,8)),
			11316 => std_logic_vector(to_unsigned( 55,8)),
			11317 => std_logic_vector(to_unsigned( 88,8)),
			11318 => std_logic_vector(to_unsigned( 36,8)),
			11319 => std_logic_vector(to_unsigned( 158,8)),
			11320 => std_logic_vector(to_unsigned( 47,8)),
			11321 => std_logic_vector(to_unsigned( 79,8)),
			11322 => std_logic_vector(to_unsigned( 50,8)),
			11323 => std_logic_vector(to_unsigned( 69,8)),
			11324 => std_logic_vector(to_unsigned( 95,8)),
			11325 => std_logic_vector(to_unsigned( 77,8)),
			11326 => std_logic_vector(to_unsigned( 176,8)),
			11327 => std_logic_vector(to_unsigned( 231,8)),
			11328 => std_logic_vector(to_unsigned( 242,8)),
			11329 => std_logic_vector(to_unsigned( 131,8)),
			11330 => std_logic_vector(to_unsigned( 220,8)),
			11331 => std_logic_vector(to_unsigned( 60,8)),
			11332 => std_logic_vector(to_unsigned( 193,8)),
			11333 => std_logic_vector(to_unsigned( 169,8)),
			11334 => std_logic_vector(to_unsigned( 63,8)),
			11335 => std_logic_vector(to_unsigned( 81,8)),
			11336 => std_logic_vector(to_unsigned( 43,8)),
			11337 => std_logic_vector(to_unsigned( 29,8)),
			11338 => std_logic_vector(to_unsigned( 147,8)),
			11339 => std_logic_vector(to_unsigned( 109,8)),
			11340 => std_logic_vector(to_unsigned( 33,8)),
			11341 => std_logic_vector(to_unsigned( 150,8)),
			11342 => std_logic_vector(to_unsigned( 10,8)),
			11343 => std_logic_vector(to_unsigned( 223,8)),
			11344 => std_logic_vector(to_unsigned( 69,8)),
			11345 => std_logic_vector(to_unsigned( 189,8)),
			11346 => std_logic_vector(to_unsigned( 84,8)),
			11347 => std_logic_vector(to_unsigned( 174,8)),
			11348 => std_logic_vector(to_unsigned( 137,8)),
			11349 => std_logic_vector(to_unsigned( 21,8)),
			11350 => std_logic_vector(to_unsigned( 23,8)),
			11351 => std_logic_vector(to_unsigned( 237,8)),
			11352 => std_logic_vector(to_unsigned( 177,8)),
			11353 => std_logic_vector(to_unsigned( 253,8)),
			11354 => std_logic_vector(to_unsigned( 17,8)),
			11355 => std_logic_vector(to_unsigned( 102,8)),
			11356 => std_logic_vector(to_unsigned( 47,8)),
			11357 => std_logic_vector(to_unsigned( 124,8)),
			11358 => std_logic_vector(to_unsigned( 202,8)),
			11359 => std_logic_vector(to_unsigned( 142,8)),
			11360 => std_logic_vector(to_unsigned( 126,8)),
			11361 => std_logic_vector(to_unsigned( 7,8)),
			11362 => std_logic_vector(to_unsigned( 152,8)),
			11363 => std_logic_vector(to_unsigned( 156,8)),
			11364 => std_logic_vector(to_unsigned( 93,8)),
			11365 => std_logic_vector(to_unsigned( 140,8)),
			11366 => std_logic_vector(to_unsigned( 78,8)),
			11367 => std_logic_vector(to_unsigned( 8,8)),
			11368 => std_logic_vector(to_unsigned( 137,8)),
			11369 => std_logic_vector(to_unsigned( 93,8)),
			11370 => std_logic_vector(to_unsigned( 114,8)),
			11371 => std_logic_vector(to_unsigned( 98,8)),
			11372 => std_logic_vector(to_unsigned( 44,8)),
			11373 => std_logic_vector(to_unsigned( 17,8)),
			11374 => std_logic_vector(to_unsigned( 66,8)),
			11375 => std_logic_vector(to_unsigned( 170,8)),
			11376 => std_logic_vector(to_unsigned( 113,8)),
			11377 => std_logic_vector(to_unsigned( 69,8)),
			11378 => std_logic_vector(to_unsigned( 230,8)),
			11379 => std_logic_vector(to_unsigned( 205,8)),
			11380 => std_logic_vector(to_unsigned( 115,8)),
			11381 => std_logic_vector(to_unsigned( 159,8)),
			11382 => std_logic_vector(to_unsigned( 15,8)),
			11383 => std_logic_vector(to_unsigned( 75,8)),
			11384 => std_logic_vector(to_unsigned( 68,8)),
			11385 => std_logic_vector(to_unsigned( 67,8)),
			11386 => std_logic_vector(to_unsigned( 59,8)),
			11387 => std_logic_vector(to_unsigned( 155,8)),
			11388 => std_logic_vector(to_unsigned( 241,8)),
			11389 => std_logic_vector(to_unsigned( 188,8)),
			11390 => std_logic_vector(to_unsigned( 148,8)),
			11391 => std_logic_vector(to_unsigned( 51,8)),
			11392 => std_logic_vector(to_unsigned( 143,8)),
			11393 => std_logic_vector(to_unsigned( 63,8)),
			11394 => std_logic_vector(to_unsigned( 141,8)),
			11395 => std_logic_vector(to_unsigned( 195,8)),
			11396 => std_logic_vector(to_unsigned( 202,8)),
			11397 => std_logic_vector(to_unsigned( 23,8)),
			11398 => std_logic_vector(to_unsigned( 1,8)),
			11399 => std_logic_vector(to_unsigned( 175,8)),
			11400 => std_logic_vector(to_unsigned( 20,8)),
			11401 => std_logic_vector(to_unsigned( 131,8)),
			11402 => std_logic_vector(to_unsigned( 109,8)),
			11403 => std_logic_vector(to_unsigned( 248,8)),
			11404 => std_logic_vector(to_unsigned( 108,8)),
			11405 => std_logic_vector(to_unsigned( 148,8)),
			11406 => std_logic_vector(to_unsigned( 57,8)),
			11407 => std_logic_vector(to_unsigned( 175,8)),
			11408 => std_logic_vector(to_unsigned( 154,8)),
			11409 => std_logic_vector(to_unsigned( 181,8)),
			11410 => std_logic_vector(to_unsigned( 235,8)),
			11411 => std_logic_vector(to_unsigned( 52,8)),
			11412 => std_logic_vector(to_unsigned( 108,8)),
			11413 => std_logic_vector(to_unsigned( 17,8)),
			11414 => std_logic_vector(to_unsigned( 14,8)),
			11415 => std_logic_vector(to_unsigned( 246,8)),
			11416 => std_logic_vector(to_unsigned( 164,8)),
			11417 => std_logic_vector(to_unsigned( 230,8)),
			11418 => std_logic_vector(to_unsigned( 139,8)),
			11419 => std_logic_vector(to_unsigned( 74,8)),
			11420 => std_logic_vector(to_unsigned( 243,8)),
			11421 => std_logic_vector(to_unsigned( 217,8)),
			11422 => std_logic_vector(to_unsigned( 103,8)),
			11423 => std_logic_vector(to_unsigned( 124,8)),
			11424 => std_logic_vector(to_unsigned( 119,8)),
			11425 => std_logic_vector(to_unsigned( 157,8)),
			11426 => std_logic_vector(to_unsigned( 50,8)),
			11427 => std_logic_vector(to_unsigned( 91,8)),
			11428 => std_logic_vector(to_unsigned( 140,8)),
			11429 => std_logic_vector(to_unsigned( 133,8)),
			11430 => std_logic_vector(to_unsigned( 57,8)),
			11431 => std_logic_vector(to_unsigned( 10,8)),
			11432 => std_logic_vector(to_unsigned( 183,8)),
			11433 => std_logic_vector(to_unsigned( 127,8)),
			11434 => std_logic_vector(to_unsigned( 7,8)),
			11435 => std_logic_vector(to_unsigned( 65,8)),
			11436 => std_logic_vector(to_unsigned( 250,8)),
			11437 => std_logic_vector(to_unsigned( 124,8)),
			11438 => std_logic_vector(to_unsigned( 45,8)),
			11439 => std_logic_vector(to_unsigned( 169,8)),
			11440 => std_logic_vector(to_unsigned( 20,8)),
			11441 => std_logic_vector(to_unsigned( 240,8)),
			11442 => std_logic_vector(to_unsigned( 7,8)),
			11443 => std_logic_vector(to_unsigned( 195,8)),
			11444 => std_logic_vector(to_unsigned( 117,8)),
			11445 => std_logic_vector(to_unsigned( 31,8)),
			11446 => std_logic_vector(to_unsigned( 19,8)),
			11447 => std_logic_vector(to_unsigned( 247,8)),
			11448 => std_logic_vector(to_unsigned( 67,8)),
			11449 => std_logic_vector(to_unsigned( 183,8)),
			11450 => std_logic_vector(to_unsigned( 89,8)),
			11451 => std_logic_vector(to_unsigned( 19,8)),
			11452 => std_logic_vector(to_unsigned( 233,8)),
			11453 => std_logic_vector(to_unsigned( 135,8)),
			11454 => std_logic_vector(to_unsigned( 247,8)),
			11455 => std_logic_vector(to_unsigned( 11,8)),
			11456 => std_logic_vector(to_unsigned( 252,8)),
			11457 => std_logic_vector(to_unsigned( 5,8)),
			11458 => std_logic_vector(to_unsigned( 68,8)),
			11459 => std_logic_vector(to_unsigned( 190,8)),
			11460 => std_logic_vector(to_unsigned( 111,8)),
			11461 => std_logic_vector(to_unsigned( 94,8)),
			11462 => std_logic_vector(to_unsigned( 201,8)),
			11463 => std_logic_vector(to_unsigned( 60,8)),
			11464 => std_logic_vector(to_unsigned( 96,8)),
			11465 => std_logic_vector(to_unsigned( 29,8)),
			11466 => std_logic_vector(to_unsigned( 20,8)),
			11467 => std_logic_vector(to_unsigned( 71,8)),
			11468 => std_logic_vector(to_unsigned( 46,8)),
			11469 => std_logic_vector(to_unsigned( 182,8)),
			11470 => std_logic_vector(to_unsigned( 154,8)),
			11471 => std_logic_vector(to_unsigned( 180,8)),
			11472 => std_logic_vector(to_unsigned( 75,8)),
			11473 => std_logic_vector(to_unsigned( 52,8)),
			11474 => std_logic_vector(to_unsigned( 75,8)),
			11475 => std_logic_vector(to_unsigned( 70,8)),
			11476 => std_logic_vector(to_unsigned( 227,8)),
			11477 => std_logic_vector(to_unsigned( 63,8)),
			11478 => std_logic_vector(to_unsigned( 41,8)),
			11479 => std_logic_vector(to_unsigned( 147,8)),
			11480 => std_logic_vector(to_unsigned( 9,8)),
			11481 => std_logic_vector(to_unsigned( 219,8)),
			11482 => std_logic_vector(to_unsigned( 137,8)),
			11483 => std_logic_vector(to_unsigned( 218,8)),
			11484 => std_logic_vector(to_unsigned( 195,8)),
			11485 => std_logic_vector(to_unsigned( 170,8)),
			11486 => std_logic_vector(to_unsigned( 127,8)),
			11487 => std_logic_vector(to_unsigned( 246,8)),
			11488 => std_logic_vector(to_unsigned( 160,8)),
			11489 => std_logic_vector(to_unsigned( 166,8)),
			11490 => std_logic_vector(to_unsigned( 75,8)),
			11491 => std_logic_vector(to_unsigned( 61,8)),
			11492 => std_logic_vector(to_unsigned( 180,8)),
			11493 => std_logic_vector(to_unsigned( 221,8)),
			11494 => std_logic_vector(to_unsigned( 194,8)),
			11495 => std_logic_vector(to_unsigned( 58,8)),
			11496 => std_logic_vector(to_unsigned( 168,8)),
			11497 => std_logic_vector(to_unsigned( 55,8)),
			11498 => std_logic_vector(to_unsigned( 124,8)),
			11499 => std_logic_vector(to_unsigned( 134,8)),
			11500 => std_logic_vector(to_unsigned( 119,8)),
			11501 => std_logic_vector(to_unsigned( 12,8)),
			11502 => std_logic_vector(to_unsigned( 92,8)),
			11503 => std_logic_vector(to_unsigned( 82,8)),
			11504 => std_logic_vector(to_unsigned( 59,8)),
			11505 => std_logic_vector(to_unsigned( 76,8)),
			11506 => std_logic_vector(to_unsigned( 198,8)),
			11507 => std_logic_vector(to_unsigned( 255,8)),
			11508 => std_logic_vector(to_unsigned( 13,8)),
			11509 => std_logic_vector(to_unsigned( 226,8)),
			11510 => std_logic_vector(to_unsigned( 216,8)),
			11511 => std_logic_vector(to_unsigned( 124,8)),
			11512 => std_logic_vector(to_unsigned( 252,8)),
			11513 => std_logic_vector(to_unsigned( 232,8)),
			11514 => std_logic_vector(to_unsigned( 6,8)),
			11515 => std_logic_vector(to_unsigned( 120,8)),
			11516 => std_logic_vector(to_unsigned( 190,8)),
			11517 => std_logic_vector(to_unsigned( 139,8)),
			11518 => std_logic_vector(to_unsigned( 31,8)),
			11519 => std_logic_vector(to_unsigned( 83,8)),
			11520 => std_logic_vector(to_unsigned( 197,8)),
			11521 => std_logic_vector(to_unsigned( 30,8)),
			11522 => std_logic_vector(to_unsigned( 50,8)),
			11523 => std_logic_vector(to_unsigned( 236,8)),
			11524 => std_logic_vector(to_unsigned( 156,8)),
			11525 => std_logic_vector(to_unsigned( 215,8)),
			11526 => std_logic_vector(to_unsigned( 170,8)),
			11527 => std_logic_vector(to_unsigned( 253,8)),
			11528 => std_logic_vector(to_unsigned( 116,8)),
			11529 => std_logic_vector(to_unsigned( 244,8)),
			11530 => std_logic_vector(to_unsigned( 187,8)),
			11531 => std_logic_vector(to_unsigned( 7,8)),
			11532 => std_logic_vector(to_unsigned( 185,8)),
			11533 => std_logic_vector(to_unsigned( 162,8)),
			11534 => std_logic_vector(to_unsigned( 38,8)),
			11535 => std_logic_vector(to_unsigned( 42,8)),
			11536 => std_logic_vector(to_unsigned( 89,8)),
			11537 => std_logic_vector(to_unsigned( 114,8)),
			11538 => std_logic_vector(to_unsigned( 154,8)),
			11539 => std_logic_vector(to_unsigned( 43,8)),
			11540 => std_logic_vector(to_unsigned( 66,8)),
			11541 => std_logic_vector(to_unsigned( 233,8)),
			11542 => std_logic_vector(to_unsigned( 77,8)),
			11543 => std_logic_vector(to_unsigned( 29,8)),
			11544 => std_logic_vector(to_unsigned( 211,8)),
			11545 => std_logic_vector(to_unsigned( 250,8)),
			11546 => std_logic_vector(to_unsigned( 145,8)),
			11547 => std_logic_vector(to_unsigned( 216,8)),
			11548 => std_logic_vector(to_unsigned( 101,8)),
			11549 => std_logic_vector(to_unsigned( 145,8)),
			11550 => std_logic_vector(to_unsigned( 179,8)),
			11551 => std_logic_vector(to_unsigned( 67,8)),
			11552 => std_logic_vector(to_unsigned( 21,8)),
			11553 => std_logic_vector(to_unsigned( 139,8)),
			11554 => std_logic_vector(to_unsigned( 208,8)),
			11555 => std_logic_vector(to_unsigned( 12,8)),
			11556 => std_logic_vector(to_unsigned( 197,8)),
			11557 => std_logic_vector(to_unsigned( 61,8)),
			11558 => std_logic_vector(to_unsigned( 142,8)),
			11559 => std_logic_vector(to_unsigned( 223,8)),
			11560 => std_logic_vector(to_unsigned( 4,8)),
			11561 => std_logic_vector(to_unsigned( 162,8)),
			11562 => std_logic_vector(to_unsigned( 181,8)),
			11563 => std_logic_vector(to_unsigned( 192,8)),
			11564 => std_logic_vector(to_unsigned( 91,8)),
			11565 => std_logic_vector(to_unsigned( 91,8)),
			11566 => std_logic_vector(to_unsigned( 151,8)),
			11567 => std_logic_vector(to_unsigned( 142,8)),
			11568 => std_logic_vector(to_unsigned( 167,8)),
			11569 => std_logic_vector(to_unsigned( 217,8)),
			11570 => std_logic_vector(to_unsigned( 183,8)),
			11571 => std_logic_vector(to_unsigned( 236,8)),
			11572 => std_logic_vector(to_unsigned( 127,8)),
			11573 => std_logic_vector(to_unsigned( 62,8)),
			11574 => std_logic_vector(to_unsigned( 228,8)),
			11575 => std_logic_vector(to_unsigned( 106,8)),
			11576 => std_logic_vector(to_unsigned( 63,8)),
			11577 => std_logic_vector(to_unsigned( 120,8)),
			11578 => std_logic_vector(to_unsigned( 245,8)),
			11579 => std_logic_vector(to_unsigned( 96,8)),
			11580 => std_logic_vector(to_unsigned( 249,8)),
			11581 => std_logic_vector(to_unsigned( 213,8)),
			11582 => std_logic_vector(to_unsigned( 77,8)),
			11583 => std_logic_vector(to_unsigned( 37,8)),
			11584 => std_logic_vector(to_unsigned( 240,8)),
			11585 => std_logic_vector(to_unsigned( 166,8)),
			11586 => std_logic_vector(to_unsigned( 41,8)),
			11587 => std_logic_vector(to_unsigned( 10,8)),
			11588 => std_logic_vector(to_unsigned( 108,8)),
			11589 => std_logic_vector(to_unsigned( 98,8)),
			11590 => std_logic_vector(to_unsigned( 125,8)),
			11591 => std_logic_vector(to_unsigned( 162,8)),
			11592 => std_logic_vector(to_unsigned( 30,8)),
			11593 => std_logic_vector(to_unsigned( 37,8)),
			11594 => std_logic_vector(to_unsigned( 36,8)),
			11595 => std_logic_vector(to_unsigned( 157,8)),
			11596 => std_logic_vector(to_unsigned( 243,8)),
			11597 => std_logic_vector(to_unsigned( 97,8)),
			11598 => std_logic_vector(to_unsigned( 161,8)),
			11599 => std_logic_vector(to_unsigned( 104,8)),
			11600 => std_logic_vector(to_unsigned( 66,8)),
			11601 => std_logic_vector(to_unsigned( 91,8)),
			11602 => std_logic_vector(to_unsigned( 175,8)),
			11603 => std_logic_vector(to_unsigned( 9,8)),
			11604 => std_logic_vector(to_unsigned( 212,8)),
			11605 => std_logic_vector(to_unsigned( 16,8)),
			11606 => std_logic_vector(to_unsigned( 250,8)),
			11607 => std_logic_vector(to_unsigned( 238,8)),
			11608 => std_logic_vector(to_unsigned( 189,8)),
			11609 => std_logic_vector(to_unsigned( 121,8)),
			11610 => std_logic_vector(to_unsigned( 74,8)),
			11611 => std_logic_vector(to_unsigned( 225,8)),
			11612 => std_logic_vector(to_unsigned( 241,8)),
			11613 => std_logic_vector(to_unsigned( 50,8)),
			11614 => std_logic_vector(to_unsigned( 219,8)),
			11615 => std_logic_vector(to_unsigned( 119,8)),
			11616 => std_logic_vector(to_unsigned( 220,8)),
			11617 => std_logic_vector(to_unsigned( 132,8)),
			11618 => std_logic_vector(to_unsigned( 126,8)),
			11619 => std_logic_vector(to_unsigned( 193,8)),
			11620 => std_logic_vector(to_unsigned( 221,8)),
			11621 => std_logic_vector(to_unsigned( 47,8)),
			11622 => std_logic_vector(to_unsigned( 136,8)),
			11623 => std_logic_vector(to_unsigned( 254,8)),
			11624 => std_logic_vector(to_unsigned( 241,8)),
			11625 => std_logic_vector(to_unsigned( 77,8)),
			11626 => std_logic_vector(to_unsigned( 186,8)),
			11627 => std_logic_vector(to_unsigned( 4,8)),
			11628 => std_logic_vector(to_unsigned( 43,8)),
			11629 => std_logic_vector(to_unsigned( 21,8)),
			11630 => std_logic_vector(to_unsigned( 111,8)),
			11631 => std_logic_vector(to_unsigned( 9,8)),
			11632 => std_logic_vector(to_unsigned( 107,8)),
			11633 => std_logic_vector(to_unsigned( 176,8)),
			11634 => std_logic_vector(to_unsigned( 244,8)),
			11635 => std_logic_vector(to_unsigned( 158,8)),
			11636 => std_logic_vector(to_unsigned( 38,8)),
			11637 => std_logic_vector(to_unsigned( 150,8)),
			11638 => std_logic_vector(to_unsigned( 234,8)),
			11639 => std_logic_vector(to_unsigned( 135,8)),
			11640 => std_logic_vector(to_unsigned( 6,8)),
			11641 => std_logic_vector(to_unsigned( 0,8)),
			11642 => std_logic_vector(to_unsigned( 154,8)),
			11643 => std_logic_vector(to_unsigned( 117,8)),
			11644 => std_logic_vector(to_unsigned( 174,8)),
			11645 => std_logic_vector(to_unsigned( 183,8)),
			11646 => std_logic_vector(to_unsigned( 239,8)),
			11647 => std_logic_vector(to_unsigned( 121,8)),
			11648 => std_logic_vector(to_unsigned( 17,8)),
			11649 => std_logic_vector(to_unsigned( 77,8)),
			11650 => std_logic_vector(to_unsigned( 235,8)),
			11651 => std_logic_vector(to_unsigned( 41,8)),
			11652 => std_logic_vector(to_unsigned( 71,8)),
			11653 => std_logic_vector(to_unsigned( 93,8)),
			11654 => std_logic_vector(to_unsigned( 179,8)),
			11655 => std_logic_vector(to_unsigned( 41,8)),
			11656 => std_logic_vector(to_unsigned( 196,8)),
			11657 => std_logic_vector(to_unsigned( 121,8)),
			11658 => std_logic_vector(to_unsigned( 125,8)),
			11659 => std_logic_vector(to_unsigned( 232,8)),
			11660 => std_logic_vector(to_unsigned( 103,8)),
			11661 => std_logic_vector(to_unsigned( 52,8)),
			11662 => std_logic_vector(to_unsigned( 121,8)),
			11663 => std_logic_vector(to_unsigned( 156,8)),
			11664 => std_logic_vector(to_unsigned( 195,8)),
			11665 => std_logic_vector(to_unsigned( 200,8)),
			11666 => std_logic_vector(to_unsigned( 220,8)),
			11667 => std_logic_vector(to_unsigned( 120,8)),
			11668 => std_logic_vector(to_unsigned( 246,8)),
			11669 => std_logic_vector(to_unsigned( 116,8)),
			11670 => std_logic_vector(to_unsigned( 9,8)),
			11671 => std_logic_vector(to_unsigned( 21,8)),
			11672 => std_logic_vector(to_unsigned( 23,8)),
			11673 => std_logic_vector(to_unsigned( 253,8)),
			11674 => std_logic_vector(to_unsigned( 60,8)),
			11675 => std_logic_vector(to_unsigned( 119,8)),
			11676 => std_logic_vector(to_unsigned( 189,8)),
			11677 => std_logic_vector(to_unsigned( 195,8)),
			11678 => std_logic_vector(to_unsigned( 247,8)),
			11679 => std_logic_vector(to_unsigned( 226,8)),
			11680 => std_logic_vector(to_unsigned( 50,8)),
			11681 => std_logic_vector(to_unsigned( 106,8)),
			11682 => std_logic_vector(to_unsigned( 86,8)),
			11683 => std_logic_vector(to_unsigned( 147,8)),
			11684 => std_logic_vector(to_unsigned( 8,8)),
			11685 => std_logic_vector(to_unsigned( 252,8)),
			11686 => std_logic_vector(to_unsigned( 217,8)),
			11687 => std_logic_vector(to_unsigned( 209,8)),
			11688 => std_logic_vector(to_unsigned( 22,8)),
			11689 => std_logic_vector(to_unsigned( 254,8)),
			11690 => std_logic_vector(to_unsigned( 191,8)),
			11691 => std_logic_vector(to_unsigned( 234,8)),
			11692 => std_logic_vector(to_unsigned( 4,8)),
			11693 => std_logic_vector(to_unsigned( 51,8)),
			11694 => std_logic_vector(to_unsigned( 139,8)),
			11695 => std_logic_vector(to_unsigned( 140,8)),
			11696 => std_logic_vector(to_unsigned( 14,8)),
			11697 => std_logic_vector(to_unsigned( 221,8)),
			11698 => std_logic_vector(to_unsigned( 129,8)),
			11699 => std_logic_vector(to_unsigned( 131,8)),
			11700 => std_logic_vector(to_unsigned( 177,8)),
			11701 => std_logic_vector(to_unsigned( 225,8)),
			11702 => std_logic_vector(to_unsigned( 87,8)),
			11703 => std_logic_vector(to_unsigned( 5,8)),
			11704 => std_logic_vector(to_unsigned( 168,8)),
			11705 => std_logic_vector(to_unsigned( 14,8)),
			11706 => std_logic_vector(to_unsigned( 53,8)),
			11707 => std_logic_vector(to_unsigned( 150,8)),
			11708 => std_logic_vector(to_unsigned( 235,8)),
			11709 => std_logic_vector(to_unsigned( 214,8)),
			11710 => std_logic_vector(to_unsigned( 91,8)),
			11711 => std_logic_vector(to_unsigned( 15,8)),
			11712 => std_logic_vector(to_unsigned( 109,8)),
			11713 => std_logic_vector(to_unsigned( 99,8)),
			11714 => std_logic_vector(to_unsigned( 179,8)),
			11715 => std_logic_vector(to_unsigned( 28,8)),
			11716 => std_logic_vector(to_unsigned( 102,8)),
			11717 => std_logic_vector(to_unsigned( 126,8)),
			11718 => std_logic_vector(to_unsigned( 213,8)),
			11719 => std_logic_vector(to_unsigned( 92,8)),
			11720 => std_logic_vector(to_unsigned( 4,8)),
			11721 => std_logic_vector(to_unsigned( 230,8)),
			11722 => std_logic_vector(to_unsigned( 65,8)),
			11723 => std_logic_vector(to_unsigned( 3,8)),
			11724 => std_logic_vector(to_unsigned( 139,8)),
			11725 => std_logic_vector(to_unsigned( 32,8)),
			11726 => std_logic_vector(to_unsigned( 44,8)),
			11727 => std_logic_vector(to_unsigned( 17,8)),
			11728 => std_logic_vector(to_unsigned( 31,8)),
			11729 => std_logic_vector(to_unsigned( 49,8)),
			11730 => std_logic_vector(to_unsigned( 187,8)),
			11731 => std_logic_vector(to_unsigned( 236,8)),
			11732 => std_logic_vector(to_unsigned( 26,8)),
			11733 => std_logic_vector(to_unsigned( 53,8)),
			11734 => std_logic_vector(to_unsigned( 240,8)),
			11735 => std_logic_vector(to_unsigned( 37,8)),
			11736 => std_logic_vector(to_unsigned( 96,8)),
			11737 => std_logic_vector(to_unsigned( 221,8)),
			11738 => std_logic_vector(to_unsigned( 196,8)),
			11739 => std_logic_vector(to_unsigned( 1,8)),
			11740 => std_logic_vector(to_unsigned( 234,8)),
			11741 => std_logic_vector(to_unsigned( 173,8)),
			11742 => std_logic_vector(to_unsigned( 94,8)),
			11743 => std_logic_vector(to_unsigned( 116,8)),
			11744 => std_logic_vector(to_unsigned( 203,8)),
			11745 => std_logic_vector(to_unsigned( 96,8)),
			11746 => std_logic_vector(to_unsigned( 30,8)),
			11747 => std_logic_vector(to_unsigned( 211,8)),
			11748 => std_logic_vector(to_unsigned( 163,8)),
			11749 => std_logic_vector(to_unsigned( 77,8)),
			11750 => std_logic_vector(to_unsigned( 44,8)),
			11751 => std_logic_vector(to_unsigned( 142,8)),
			11752 => std_logic_vector(to_unsigned( 154,8)),
			11753 => std_logic_vector(to_unsigned( 124,8)),
			11754 => std_logic_vector(to_unsigned( 238,8)),
			11755 => std_logic_vector(to_unsigned( 87,8)),
			11756 => std_logic_vector(to_unsigned( 49,8)),
			11757 => std_logic_vector(to_unsigned( 6,8)),
			11758 => std_logic_vector(to_unsigned( 204,8)),
			11759 => std_logic_vector(to_unsigned( 197,8)),
			11760 => std_logic_vector(to_unsigned( 187,8)),
			11761 => std_logic_vector(to_unsigned( 201,8)),
			11762 => std_logic_vector(to_unsigned( 41,8)),
			11763 => std_logic_vector(to_unsigned( 130,8)),
			11764 => std_logic_vector(to_unsigned( 12,8)),
			11765 => std_logic_vector(to_unsigned( 159,8)),
			11766 => std_logic_vector(to_unsigned( 9,8)),
			11767 => std_logic_vector(to_unsigned( 231,8)),
			11768 => std_logic_vector(to_unsigned( 153,8)),
			11769 => std_logic_vector(to_unsigned( 120,8)),
			11770 => std_logic_vector(to_unsigned( 136,8)),
			11771 => std_logic_vector(to_unsigned( 220,8)),
			11772 => std_logic_vector(to_unsigned( 25,8)),
			11773 => std_logic_vector(to_unsigned( 248,8)),
			11774 => std_logic_vector(to_unsigned( 21,8)),
			11775 => std_logic_vector(to_unsigned( 176,8)),
			11776 => std_logic_vector(to_unsigned( 154,8)),
			11777 => std_logic_vector(to_unsigned( 154,8)),
			11778 => std_logic_vector(to_unsigned( 189,8)),
			11779 => std_logic_vector(to_unsigned( 100,8)),
			11780 => std_logic_vector(to_unsigned( 17,8)),
			11781 => std_logic_vector(to_unsigned( 119,8)),
			11782 => std_logic_vector(to_unsigned( 6,8)),
			11783 => std_logic_vector(to_unsigned( 122,8)),
			11784 => std_logic_vector(to_unsigned( 204,8)),
			11785 => std_logic_vector(to_unsigned( 226,8)),
			11786 => std_logic_vector(to_unsigned( 180,8)),
			11787 => std_logic_vector(to_unsigned( 242,8)),
			11788 => std_logic_vector(to_unsigned( 72,8)),
			11789 => std_logic_vector(to_unsigned( 246,8)),
			11790 => std_logic_vector(to_unsigned( 27,8)),
			11791 => std_logic_vector(to_unsigned( 98,8)),
			11792 => std_logic_vector(to_unsigned( 231,8)),
			11793 => std_logic_vector(to_unsigned( 70,8)),
			11794 => std_logic_vector(to_unsigned( 252,8)),
			11795 => std_logic_vector(to_unsigned( 17,8)),
			11796 => std_logic_vector(to_unsigned( 26,8)),
			11797 => std_logic_vector(to_unsigned( 216,8)),
			11798 => std_logic_vector(to_unsigned( 101,8)),
			11799 => std_logic_vector(to_unsigned( 146,8)),
			11800 => std_logic_vector(to_unsigned( 87,8)),
			11801 => std_logic_vector(to_unsigned( 6,8)),
			11802 => std_logic_vector(to_unsigned( 8,8)),
			11803 => std_logic_vector(to_unsigned( 173,8)),
			11804 => std_logic_vector(to_unsigned( 112,8)),
			11805 => std_logic_vector(to_unsigned( 21,8)),
			11806 => std_logic_vector(to_unsigned( 20,8)),
			11807 => std_logic_vector(to_unsigned( 74,8)),
			11808 => std_logic_vector(to_unsigned( 147,8)),
			11809 => std_logic_vector(to_unsigned( 42,8)),
			11810 => std_logic_vector(to_unsigned( 130,8)),
			11811 => std_logic_vector(to_unsigned( 85,8)),
			11812 => std_logic_vector(to_unsigned( 200,8)),
			11813 => std_logic_vector(to_unsigned( 113,8)),
			11814 => std_logic_vector(to_unsigned( 214,8)),
			11815 => std_logic_vector(to_unsigned( 117,8)),
			11816 => std_logic_vector(to_unsigned( 233,8)),
			11817 => std_logic_vector(to_unsigned( 237,8)),
			11818 => std_logic_vector(to_unsigned( 168,8)),
			11819 => std_logic_vector(to_unsigned( 72,8)),
			11820 => std_logic_vector(to_unsigned( 189,8)),
			11821 => std_logic_vector(to_unsigned( 186,8)),
			11822 => std_logic_vector(to_unsigned( 237,8)),
			11823 => std_logic_vector(to_unsigned( 110,8)),
			11824 => std_logic_vector(to_unsigned( 31,8)),
			11825 => std_logic_vector(to_unsigned( 20,8)),
			11826 => std_logic_vector(to_unsigned( 180,8)),
			11827 => std_logic_vector(to_unsigned( 139,8)),
			11828 => std_logic_vector(to_unsigned( 115,8)),
			11829 => std_logic_vector(to_unsigned( 243,8)),
			11830 => std_logic_vector(to_unsigned( 18,8)),
			11831 => std_logic_vector(to_unsigned( 193,8)),
			11832 => std_logic_vector(to_unsigned( 182,8)),
			11833 => std_logic_vector(to_unsigned( 143,8)),
			11834 => std_logic_vector(to_unsigned( 68,8)),
			11835 => std_logic_vector(to_unsigned( 98,8)),
			11836 => std_logic_vector(to_unsigned( 102,8)),
			11837 => std_logic_vector(to_unsigned( 174,8)),
			11838 => std_logic_vector(to_unsigned( 12,8)),
			11839 => std_logic_vector(to_unsigned( 221,8)),
			11840 => std_logic_vector(to_unsigned( 161,8)),
			11841 => std_logic_vector(to_unsigned( 107,8)),
			11842 => std_logic_vector(to_unsigned( 210,8)),
			11843 => std_logic_vector(to_unsigned( 54,8)),
			11844 => std_logic_vector(to_unsigned( 166,8)),
			11845 => std_logic_vector(to_unsigned( 165,8)),
			11846 => std_logic_vector(to_unsigned( 136,8)),
			11847 => std_logic_vector(to_unsigned( 52,8)),
			11848 => std_logic_vector(to_unsigned( 78,8)),
			11849 => std_logic_vector(to_unsigned( 239,8)),
			11850 => std_logic_vector(to_unsigned( 13,8)),
			11851 => std_logic_vector(to_unsigned( 51,8)),
			11852 => std_logic_vector(to_unsigned( 228,8)),
			11853 => std_logic_vector(to_unsigned( 105,8)),
			11854 => std_logic_vector(to_unsigned( 160,8)),
			11855 => std_logic_vector(to_unsigned( 203,8)),
			11856 => std_logic_vector(to_unsigned( 209,8)),
			11857 => std_logic_vector(to_unsigned( 106,8)),
			11858 => std_logic_vector(to_unsigned( 128,8)),
			11859 => std_logic_vector(to_unsigned( 188,8)),
			11860 => std_logic_vector(to_unsigned( 168,8)),
			11861 => std_logic_vector(to_unsigned( 214,8)),
			11862 => std_logic_vector(to_unsigned( 35,8)),
			11863 => std_logic_vector(to_unsigned( 231,8)),
			11864 => std_logic_vector(to_unsigned( 192,8)),
			11865 => std_logic_vector(to_unsigned( 83,8)),
			11866 => std_logic_vector(to_unsigned( 146,8)),
			11867 => std_logic_vector(to_unsigned( 247,8)),
			11868 => std_logic_vector(to_unsigned( 56,8)),
			11869 => std_logic_vector(to_unsigned( 158,8)),
			11870 => std_logic_vector(to_unsigned( 170,8)),
			11871 => std_logic_vector(to_unsigned( 189,8)),
			11872 => std_logic_vector(to_unsigned( 224,8)),
			11873 => std_logic_vector(to_unsigned( 209,8)),
			11874 => std_logic_vector(to_unsigned( 215,8)),
			11875 => std_logic_vector(to_unsigned( 197,8)),
			11876 => std_logic_vector(to_unsigned( 114,8)),
			11877 => std_logic_vector(to_unsigned( 20,8)),
			11878 => std_logic_vector(to_unsigned( 17,8)),
			11879 => std_logic_vector(to_unsigned( 154,8)),
			11880 => std_logic_vector(to_unsigned( 30,8)),
			11881 => std_logic_vector(to_unsigned( 5,8)),
			11882 => std_logic_vector(to_unsigned( 118,8)),
			11883 => std_logic_vector(to_unsigned( 38,8)),
			11884 => std_logic_vector(to_unsigned( 64,8)),
			11885 => std_logic_vector(to_unsigned( 163,8)),
			11886 => std_logic_vector(to_unsigned( 117,8)),
			11887 => std_logic_vector(to_unsigned( 5,8)),
			11888 => std_logic_vector(to_unsigned( 163,8)),
			11889 => std_logic_vector(to_unsigned( 234,8)),
			11890 => std_logic_vector(to_unsigned( 236,8)),
			11891 => std_logic_vector(to_unsigned( 202,8)),
			11892 => std_logic_vector(to_unsigned( 23,8)),
			11893 => std_logic_vector(to_unsigned( 137,8)),
			11894 => std_logic_vector(to_unsigned( 29,8)),
			11895 => std_logic_vector(to_unsigned( 98,8)),
			11896 => std_logic_vector(to_unsigned( 94,8)),
			11897 => std_logic_vector(to_unsigned( 8,8)),
			11898 => std_logic_vector(to_unsigned( 142,8)),
			11899 => std_logic_vector(to_unsigned( 175,8)),
			11900 => std_logic_vector(to_unsigned( 182,8)),
			11901 => std_logic_vector(to_unsigned( 144,8)),
			11902 => std_logic_vector(to_unsigned( 115,8)),
			11903 => std_logic_vector(to_unsigned( 45,8)),
			11904 => std_logic_vector(to_unsigned( 141,8)),
			11905 => std_logic_vector(to_unsigned( 248,8)),
			11906 => std_logic_vector(to_unsigned( 154,8)),
			11907 => std_logic_vector(to_unsigned( 104,8)),
			11908 => std_logic_vector(to_unsigned( 231,8)),
			11909 => std_logic_vector(to_unsigned( 78,8)),
			11910 => std_logic_vector(to_unsigned( 113,8)),
			11911 => std_logic_vector(to_unsigned( 44,8)),
			11912 => std_logic_vector(to_unsigned( 123,8)),
			11913 => std_logic_vector(to_unsigned( 168,8)),
			11914 => std_logic_vector(to_unsigned( 168,8)),
			11915 => std_logic_vector(to_unsigned( 156,8)),
			11916 => std_logic_vector(to_unsigned( 52,8)),
			11917 => std_logic_vector(to_unsigned( 145,8)),
			11918 => std_logic_vector(to_unsigned( 224,8)),
			11919 => std_logic_vector(to_unsigned( 212,8)),
			11920 => std_logic_vector(to_unsigned( 237,8)),
			11921 => std_logic_vector(to_unsigned( 6,8)),
			11922 => std_logic_vector(to_unsigned( 0,8)),
			11923 => std_logic_vector(to_unsigned( 174,8)),
			11924 => std_logic_vector(to_unsigned( 69,8)),
			11925 => std_logic_vector(to_unsigned( 57,8)),
			11926 => std_logic_vector(to_unsigned( 57,8)),
			11927 => std_logic_vector(to_unsigned( 54,8)),
			11928 => std_logic_vector(to_unsigned( 71,8)),
			11929 => std_logic_vector(to_unsigned( 220,8)),
			11930 => std_logic_vector(to_unsigned( 67,8)),
			11931 => std_logic_vector(to_unsigned( 198,8)),
			11932 => std_logic_vector(to_unsigned( 250,8)),
			11933 => std_logic_vector(to_unsigned( 89,8)),
			11934 => std_logic_vector(to_unsigned( 219,8)),
			11935 => std_logic_vector(to_unsigned( 96,8)),
			11936 => std_logic_vector(to_unsigned( 102,8)),
			11937 => std_logic_vector(to_unsigned( 77,8)),
			11938 => std_logic_vector(to_unsigned( 60,8)),
			11939 => std_logic_vector(to_unsigned( 145,8)),
			11940 => std_logic_vector(to_unsigned( 87,8)),
			11941 => std_logic_vector(to_unsigned( 165,8)),
			11942 => std_logic_vector(to_unsigned( 82,8)),
			11943 => std_logic_vector(to_unsigned( 158,8)),
			11944 => std_logic_vector(to_unsigned( 92,8)),
			11945 => std_logic_vector(to_unsigned( 138,8)),
			11946 => std_logic_vector(to_unsigned( 169,8)),
			11947 => std_logic_vector(to_unsigned( 95,8)),
			11948 => std_logic_vector(to_unsigned( 83,8)),
			11949 => std_logic_vector(to_unsigned( 156,8)),
			11950 => std_logic_vector(to_unsigned( 29,8)),
			11951 => std_logic_vector(to_unsigned( 26,8)),
			11952 => std_logic_vector(to_unsigned( 102,8)),
			11953 => std_logic_vector(to_unsigned( 62,8)),
			11954 => std_logic_vector(to_unsigned( 87,8)),
			11955 => std_logic_vector(to_unsigned( 80,8)),
			11956 => std_logic_vector(to_unsigned( 170,8)),
			11957 => std_logic_vector(to_unsigned( 36,8)),
			11958 => std_logic_vector(to_unsigned( 23,8)),
			11959 => std_logic_vector(to_unsigned( 101,8)),
			11960 => std_logic_vector(to_unsigned( 75,8)),
			11961 => std_logic_vector(to_unsigned( 28,8)),
			11962 => std_logic_vector(to_unsigned( 56,8)),
			11963 => std_logic_vector(to_unsigned( 187,8)),
			11964 => std_logic_vector(to_unsigned( 40,8)),
			11965 => std_logic_vector(to_unsigned( 247,8)),
			11966 => std_logic_vector(to_unsigned( 198,8)),
			11967 => std_logic_vector(to_unsigned( 22,8)),
			11968 => std_logic_vector(to_unsigned( 245,8)),
			11969 => std_logic_vector(to_unsigned( 247,8)),
			11970 => std_logic_vector(to_unsigned( 232,8)),
			11971 => std_logic_vector(to_unsigned( 176,8)),
			11972 => std_logic_vector(to_unsigned( 92,8)),
			11973 => std_logic_vector(to_unsigned( 50,8)),
			11974 => std_logic_vector(to_unsigned( 114,8)),
			11975 => std_logic_vector(to_unsigned( 170,8)),
			11976 => std_logic_vector(to_unsigned( 139,8)),
			11977 => std_logic_vector(to_unsigned( 179,8)),
			11978 => std_logic_vector(to_unsigned( 160,8)),
			11979 => std_logic_vector(to_unsigned( 107,8)),
			11980 => std_logic_vector(to_unsigned( 138,8)),
			11981 => std_logic_vector(to_unsigned( 33,8)),
			11982 => std_logic_vector(to_unsigned( 141,8)),
			11983 => std_logic_vector(to_unsigned( 123,8)),
			11984 => std_logic_vector(to_unsigned( 162,8)),
			11985 => std_logic_vector(to_unsigned( 176,8)),
			11986 => std_logic_vector(to_unsigned( 46,8)),
			11987 => std_logic_vector(to_unsigned( 128,8)),
			11988 => std_logic_vector(to_unsigned( 179,8)),
			11989 => std_logic_vector(to_unsigned( 109,8)),
			11990 => std_logic_vector(to_unsigned( 67,8)),
			11991 => std_logic_vector(to_unsigned( 92,8)),
			11992 => std_logic_vector(to_unsigned( 41,8)),
			11993 => std_logic_vector(to_unsigned( 59,8)),
			11994 => std_logic_vector(to_unsigned( 48,8)),
			11995 => std_logic_vector(to_unsigned( 131,8)),
			11996 => std_logic_vector(to_unsigned( 162,8)),
			11997 => std_logic_vector(to_unsigned( 110,8)),
			11998 => std_logic_vector(to_unsigned( 187,8)),
			11999 => std_logic_vector(to_unsigned( 39,8)),
			12000 => std_logic_vector(to_unsigned( 205,8)),
			12001 => std_logic_vector(to_unsigned( 198,8)),
			12002 => std_logic_vector(to_unsigned( 227,8)),
			12003 => std_logic_vector(to_unsigned( 121,8)),
			12004 => std_logic_vector(to_unsigned( 187,8)),
			12005 => std_logic_vector(to_unsigned( 118,8)),
			12006 => std_logic_vector(to_unsigned( 4,8)),
			12007 => std_logic_vector(to_unsigned( 171,8)),
			12008 => std_logic_vector(to_unsigned( 148,8)),
			12009 => std_logic_vector(to_unsigned( 150,8)),
			12010 => std_logic_vector(to_unsigned( 176,8)),
			12011 => std_logic_vector(to_unsigned( 20,8)),
			12012 => std_logic_vector(to_unsigned( 232,8)),
			12013 => std_logic_vector(to_unsigned( 100,8)),
			12014 => std_logic_vector(to_unsigned( 176,8)),
			12015 => std_logic_vector(to_unsigned( 186,8)),
			12016 => std_logic_vector(to_unsigned( 14,8)),
			12017 => std_logic_vector(to_unsigned( 236,8)),
			12018 => std_logic_vector(to_unsigned( 60,8)),
			12019 => std_logic_vector(to_unsigned( 135,8)),
			12020 => std_logic_vector(to_unsigned( 34,8)),
			12021 => std_logic_vector(to_unsigned( 2,8)),
			12022 => std_logic_vector(to_unsigned( 249,8)),
			12023 => std_logic_vector(to_unsigned( 241,8)),
			12024 => std_logic_vector(to_unsigned( 129,8)),
			12025 => std_logic_vector(to_unsigned( 65,8)),
			12026 => std_logic_vector(to_unsigned( 138,8)),
			12027 => std_logic_vector(to_unsigned( 101,8)),
			12028 => std_logic_vector(to_unsigned( 144,8)),
			12029 => std_logic_vector(to_unsigned( 42,8)),
			12030 => std_logic_vector(to_unsigned( 197,8)),
			12031 => std_logic_vector(to_unsigned( 228,8)),
			12032 => std_logic_vector(to_unsigned( 153,8)),
			12033 => std_logic_vector(to_unsigned( 34,8)),
			12034 => std_logic_vector(to_unsigned( 158,8)),
			12035 => std_logic_vector(to_unsigned( 174,8)),
			12036 => std_logic_vector(to_unsigned( 115,8)),
			12037 => std_logic_vector(to_unsigned( 211,8)),
			12038 => std_logic_vector(to_unsigned( 166,8)),
			12039 => std_logic_vector(to_unsigned( 19,8)),
			12040 => std_logic_vector(to_unsigned( 255,8)),
			12041 => std_logic_vector(to_unsigned( 112,8)),
			12042 => std_logic_vector(to_unsigned( 91,8)),
			12043 => std_logic_vector(to_unsigned( 30,8)),
			12044 => std_logic_vector(to_unsigned( 71,8)),
			12045 => std_logic_vector(to_unsigned( 93,8)),
			12046 => std_logic_vector(to_unsigned( 239,8)),
			12047 => std_logic_vector(to_unsigned( 114,8)),
			12048 => std_logic_vector(to_unsigned( 162,8)),
			12049 => std_logic_vector(to_unsigned( 86,8)),
			12050 => std_logic_vector(to_unsigned( 225,8)),
			12051 => std_logic_vector(to_unsigned( 125,8)),
			12052 => std_logic_vector(to_unsigned( 190,8)),
			12053 => std_logic_vector(to_unsigned( 227,8)),
			12054 => std_logic_vector(to_unsigned( 253,8)),
			12055 => std_logic_vector(to_unsigned( 167,8)),
			12056 => std_logic_vector(to_unsigned( 41,8)),
			12057 => std_logic_vector(to_unsigned( 31,8)),
			12058 => std_logic_vector(to_unsigned( 117,8)),
			12059 => std_logic_vector(to_unsigned( 37,8)),
			12060 => std_logic_vector(to_unsigned( 40,8)),
			12061 => std_logic_vector(to_unsigned( 18,8)),
			12062 => std_logic_vector(to_unsigned( 71,8)),
			12063 => std_logic_vector(to_unsigned( 99,8)),
			12064 => std_logic_vector(to_unsigned( 73,8)),
			12065 => std_logic_vector(to_unsigned( 123,8)),
			12066 => std_logic_vector(to_unsigned( 92,8)),
			12067 => std_logic_vector(to_unsigned( 173,8)),
			12068 => std_logic_vector(to_unsigned( 16,8)),
			12069 => std_logic_vector(to_unsigned( 114,8)),
			12070 => std_logic_vector(to_unsigned( 43,8)),
			12071 => std_logic_vector(to_unsigned( 116,8)),
			12072 => std_logic_vector(to_unsigned( 115,8)),
			12073 => std_logic_vector(to_unsigned( 234,8)),
			12074 => std_logic_vector(to_unsigned( 123,8)),
			12075 => std_logic_vector(to_unsigned( 163,8)),
			12076 => std_logic_vector(to_unsigned( 113,8)),
			12077 => std_logic_vector(to_unsigned( 247,8)),
			12078 => std_logic_vector(to_unsigned( 107,8)),
			12079 => std_logic_vector(to_unsigned( 99,8)),
			12080 => std_logic_vector(to_unsigned( 63,8)),
			12081 => std_logic_vector(to_unsigned( 30,8)),
			12082 => std_logic_vector(to_unsigned( 86,8)),
			12083 => std_logic_vector(to_unsigned( 82,8)),
			12084 => std_logic_vector(to_unsigned( 120,8)),
			12085 => std_logic_vector(to_unsigned( 103,8)),
			12086 => std_logic_vector(to_unsigned( 41,8)),
			12087 => std_logic_vector(to_unsigned( 192,8)),
			12088 => std_logic_vector(to_unsigned( 16,8)),
			12089 => std_logic_vector(to_unsigned( 24,8)),
			12090 => std_logic_vector(to_unsigned( 171,8)),
			12091 => std_logic_vector(to_unsigned( 187,8)),
			12092 => std_logic_vector(to_unsigned( 246,8)),
			12093 => std_logic_vector(to_unsigned( 16,8)),
			12094 => std_logic_vector(to_unsigned( 48,8)),
			12095 => std_logic_vector(to_unsigned( 228,8)),
			12096 => std_logic_vector(to_unsigned( 52,8)),
			12097 => std_logic_vector(to_unsigned( 177,8)),
			12098 => std_logic_vector(to_unsigned( 125,8)),
			12099 => std_logic_vector(to_unsigned( 221,8)),
			12100 => std_logic_vector(to_unsigned( 58,8)),
			12101 => std_logic_vector(to_unsigned( 149,8)),
			12102 => std_logic_vector(to_unsigned( 119,8)),
			12103 => std_logic_vector(to_unsigned( 242,8)),
			12104 => std_logic_vector(to_unsigned( 215,8)),
			12105 => std_logic_vector(to_unsigned( 118,8)),
			12106 => std_logic_vector(to_unsigned( 144,8)),
			12107 => std_logic_vector(to_unsigned( 141,8)),
			12108 => std_logic_vector(to_unsigned( 36,8)),
			12109 => std_logic_vector(to_unsigned( 50,8)),
			12110 => std_logic_vector(to_unsigned( 223,8)),
			12111 => std_logic_vector(to_unsigned( 99,8)),
			12112 => std_logic_vector(to_unsigned( 36,8)),
			12113 => std_logic_vector(to_unsigned( 25,8)),
			12114 => std_logic_vector(to_unsigned( 236,8)),
			12115 => std_logic_vector(to_unsigned( 176,8)),
			12116 => std_logic_vector(to_unsigned( 71,8)),
			12117 => std_logic_vector(to_unsigned( 30,8)),
			12118 => std_logic_vector(to_unsigned( 98,8)),
			12119 => std_logic_vector(to_unsigned( 150,8)),
			12120 => std_logic_vector(to_unsigned( 156,8)),
			12121 => std_logic_vector(to_unsigned( 190,8)),
			12122 => std_logic_vector(to_unsigned( 233,8)),
			12123 => std_logic_vector(to_unsigned( 219,8)),
			12124 => std_logic_vector(to_unsigned( 227,8)),
			12125 => std_logic_vector(to_unsigned( 10,8)),
			12126 => std_logic_vector(to_unsigned( 233,8)),
			12127 => std_logic_vector(to_unsigned( 142,8)),
			12128 => std_logic_vector(to_unsigned( 254,8)),
			12129 => std_logic_vector(to_unsigned( 182,8)),
			12130 => std_logic_vector(to_unsigned( 243,8)),
			12131 => std_logic_vector(to_unsigned( 154,8)),
			12132 => std_logic_vector(to_unsigned( 227,8)),
			12133 => std_logic_vector(to_unsigned( 125,8)),
			12134 => std_logic_vector(to_unsigned( 71,8)),
			12135 => std_logic_vector(to_unsigned( 112,8)),
			12136 => std_logic_vector(to_unsigned( 240,8)),
			12137 => std_logic_vector(to_unsigned( 42,8)),
			12138 => std_logic_vector(to_unsigned( 173,8)),
			12139 => std_logic_vector(to_unsigned( 108,8)),
			12140 => std_logic_vector(to_unsigned( 149,8)),
			12141 => std_logic_vector(to_unsigned( 93,8)),
			12142 => std_logic_vector(to_unsigned( 118,8)),
			12143 => std_logic_vector(to_unsigned( 35,8)),
			12144 => std_logic_vector(to_unsigned( 231,8)),
			12145 => std_logic_vector(to_unsigned( 209,8)),
			12146 => std_logic_vector(to_unsigned( 162,8)),
			12147 => std_logic_vector(to_unsigned( 196,8)),
			12148 => std_logic_vector(to_unsigned( 47,8)),
			12149 => std_logic_vector(to_unsigned( 219,8)),
			12150 => std_logic_vector(to_unsigned( 133,8)),
			12151 => std_logic_vector(to_unsigned( 3,8)),
			12152 => std_logic_vector(to_unsigned( 28,8)),
			12153 => std_logic_vector(to_unsigned( 77,8)),
			12154 => std_logic_vector(to_unsigned( 244,8)),
			12155 => std_logic_vector(to_unsigned( 71,8)),
			12156 => std_logic_vector(to_unsigned( 87,8)),
			12157 => std_logic_vector(to_unsigned( 179,8)),
			12158 => std_logic_vector(to_unsigned( 27,8)),
			12159 => std_logic_vector(to_unsigned( 235,8)),
			12160 => std_logic_vector(to_unsigned( 34,8)),
			12161 => std_logic_vector(to_unsigned( 138,8)),
			12162 => std_logic_vector(to_unsigned( 63,8)),
			12163 => std_logic_vector(to_unsigned( 98,8)),
			12164 => std_logic_vector(to_unsigned( 175,8)),
			12165 => std_logic_vector(to_unsigned( 8,8)),
			12166 => std_logic_vector(to_unsigned( 124,8)),
			12167 => std_logic_vector(to_unsigned( 143,8)),
			12168 => std_logic_vector(to_unsigned( 167,8)),
			12169 => std_logic_vector(to_unsigned( 4,8)),
			12170 => std_logic_vector(to_unsigned( 210,8)),
			12171 => std_logic_vector(to_unsigned( 36,8)),
			12172 => std_logic_vector(to_unsigned( 245,8)),
			12173 => std_logic_vector(to_unsigned( 228,8)),
			12174 => std_logic_vector(to_unsigned( 54,8)),
			12175 => std_logic_vector(to_unsigned( 157,8)),
			12176 => std_logic_vector(to_unsigned( 125,8)),
			12177 => std_logic_vector(to_unsigned( 84,8)),
			12178 => std_logic_vector(to_unsigned( 12,8)),
			12179 => std_logic_vector(to_unsigned( 214,8)),
			12180 => std_logic_vector(to_unsigned( 116,8)),
			12181 => std_logic_vector(to_unsigned( 119,8)),
			12182 => std_logic_vector(to_unsigned( 59,8)),
			12183 => std_logic_vector(to_unsigned( 72,8)),
			12184 => std_logic_vector(to_unsigned( 138,8)),
			12185 => std_logic_vector(to_unsigned( 159,8)),
			12186 => std_logic_vector(to_unsigned( 108,8)),
			12187 => std_logic_vector(to_unsigned( 226,8)),
			12188 => std_logic_vector(to_unsigned( 167,8)),
			12189 => std_logic_vector(to_unsigned( 241,8)),
			12190 => std_logic_vector(to_unsigned( 76,8)),
			12191 => std_logic_vector(to_unsigned( 172,8)),
			12192 => std_logic_vector(to_unsigned( 121,8)),
			12193 => std_logic_vector(to_unsigned( 54,8)),
			12194 => std_logic_vector(to_unsigned( 2,8)),
			12195 => std_logic_vector(to_unsigned( 183,8)),
			12196 => std_logic_vector(to_unsigned( 130,8)),
			12197 => std_logic_vector(to_unsigned( 213,8)),
			12198 => std_logic_vector(to_unsigned( 1,8)),
			12199 => std_logic_vector(to_unsigned( 127,8)),
			12200 => std_logic_vector(to_unsigned( 65,8)),
			12201 => std_logic_vector(to_unsigned( 194,8)),
			12202 => std_logic_vector(to_unsigned( 169,8)),
			12203 => std_logic_vector(to_unsigned( 78,8)),
			12204 => std_logic_vector(to_unsigned( 230,8)),
			12205 => std_logic_vector(to_unsigned( 98,8)),
			12206 => std_logic_vector(to_unsigned( 227,8)),
			12207 => std_logic_vector(to_unsigned( 114,8)),
			12208 => std_logic_vector(to_unsigned( 32,8)),
			12209 => std_logic_vector(to_unsigned( 212,8)),
			12210 => std_logic_vector(to_unsigned( 18,8)),
			12211 => std_logic_vector(to_unsigned( 25,8)),
			12212 => std_logic_vector(to_unsigned( 234,8)),
			12213 => std_logic_vector(to_unsigned( 21,8)),
			12214 => std_logic_vector(to_unsigned( 223,8)),
			12215 => std_logic_vector(to_unsigned( 59,8)),
			12216 => std_logic_vector(to_unsigned( 18,8)),
			12217 => std_logic_vector(to_unsigned( 151,8)),
			12218 => std_logic_vector(to_unsigned( 175,8)),
			12219 => std_logic_vector(to_unsigned( 124,8)),
			12220 => std_logic_vector(to_unsigned( 51,8)),
			12221 => std_logic_vector(to_unsigned( 40,8)),
			12222 => std_logic_vector(to_unsigned( 157,8)),
			12223 => std_logic_vector(to_unsigned( 109,8)),
			12224 => std_logic_vector(to_unsigned( 141,8)),
			12225 => std_logic_vector(to_unsigned( 64,8)),
			12226 => std_logic_vector(to_unsigned( 188,8)),
			12227 => std_logic_vector(to_unsigned( 132,8)),
			12228 => std_logic_vector(to_unsigned( 248,8)),
			12229 => std_logic_vector(to_unsigned( 28,8)),
			12230 => std_logic_vector(to_unsigned( 223,8)),
			12231 => std_logic_vector(to_unsigned( 75,8)),
			12232 => std_logic_vector(to_unsigned( 143,8)),
			12233 => std_logic_vector(to_unsigned( 190,8)),
			12234 => std_logic_vector(to_unsigned( 242,8)),
			12235 => std_logic_vector(to_unsigned( 102,8)),
			12236 => std_logic_vector(to_unsigned( 176,8)),
			12237 => std_logic_vector(to_unsigned( 111,8)),
			12238 => std_logic_vector(to_unsigned( 122,8)),
			12239 => std_logic_vector(to_unsigned( 219,8)),
			12240 => std_logic_vector(to_unsigned( 102,8)),
			12241 => std_logic_vector(to_unsigned( 178,8)),
			12242 => std_logic_vector(to_unsigned( 167,8)),
			12243 => std_logic_vector(to_unsigned( 224,8)),
			12244 => std_logic_vector(to_unsigned( 178,8)),
			12245 => std_logic_vector(to_unsigned( 68,8)),
			12246 => std_logic_vector(to_unsigned( 225,8)),
			12247 => std_logic_vector(to_unsigned( 199,8)),
			12248 => std_logic_vector(to_unsigned( 8,8)),
			12249 => std_logic_vector(to_unsigned( 44,8)),
			12250 => std_logic_vector(to_unsigned( 28,8)),
			12251 => std_logic_vector(to_unsigned( 173,8)),
			12252 => std_logic_vector(to_unsigned( 80,8)),
			12253 => std_logic_vector(to_unsigned( 35,8)),
			12254 => std_logic_vector(to_unsigned( 95,8)),
			12255 => std_logic_vector(to_unsigned( 209,8)),
			12256 => std_logic_vector(to_unsigned( 164,8)),
			12257 => std_logic_vector(to_unsigned( 175,8)),
			12258 => std_logic_vector(to_unsigned( 57,8)),
			12259 => std_logic_vector(to_unsigned( 103,8)),
			12260 => std_logic_vector(to_unsigned( 6,8)),
			12261 => std_logic_vector(to_unsigned( 247,8)),
			12262 => std_logic_vector(to_unsigned( 254,8)),
			12263 => std_logic_vector(to_unsigned( 72,8)),
			12264 => std_logic_vector(to_unsigned( 46,8)),
			12265 => std_logic_vector(to_unsigned( 157,8)),
			12266 => std_logic_vector(to_unsigned( 92,8)),
			12267 => std_logic_vector(to_unsigned( 61,8)),
			12268 => std_logic_vector(to_unsigned( 143,8)),
			12269 => std_logic_vector(to_unsigned( 100,8)),
			12270 => std_logic_vector(to_unsigned( 21,8)),
			12271 => std_logic_vector(to_unsigned( 139,8)),
			12272 => std_logic_vector(to_unsigned( 108,8)),
			12273 => std_logic_vector(to_unsigned( 113,8)),
			12274 => std_logic_vector(to_unsigned( 183,8)),
			12275 => std_logic_vector(to_unsigned( 191,8)),
			12276 => std_logic_vector(to_unsigned( 226,8)),
			12277 => std_logic_vector(to_unsigned( 122,8)),
			12278 => std_logic_vector(to_unsigned( 106,8)),
			12279 => std_logic_vector(to_unsigned( 174,8)),
			12280 => std_logic_vector(to_unsigned( 20,8)),
			12281 => std_logic_vector(to_unsigned( 99,8)),
			12282 => std_logic_vector(to_unsigned( 4,8)),
			12283 => std_logic_vector(to_unsigned( 214,8)),
			12284 => std_logic_vector(to_unsigned( 131,8)),
			12285 => std_logic_vector(to_unsigned( 82,8)),
			12286 => std_logic_vector(to_unsigned( 182,8)),
			12287 => std_logic_vector(to_unsigned( 23,8)),
			12288 => std_logic_vector(to_unsigned( 161,8)),
			12289 => std_logic_vector(to_unsigned( 40,8)),
			12290 => std_logic_vector(to_unsigned( 24,8)),
			12291 => std_logic_vector(to_unsigned( 59,8)),
			12292 => std_logic_vector(to_unsigned( 188,8)),
			12293 => std_logic_vector(to_unsigned( 50,8)),
			12294 => std_logic_vector(to_unsigned( 181,8)),
			12295 => std_logic_vector(to_unsigned( 232,8)),
			12296 => std_logic_vector(to_unsigned( 165,8)),
			12297 => std_logic_vector(to_unsigned( 164,8)),
			12298 => std_logic_vector(to_unsigned( 226,8)),
			12299 => std_logic_vector(to_unsigned( 207,8)),
			12300 => std_logic_vector(to_unsigned( 69,8)),
			12301 => std_logic_vector(to_unsigned( 39,8)),
			12302 => std_logic_vector(to_unsigned( 81,8)),
			12303 => std_logic_vector(to_unsigned( 251,8)),
			12304 => std_logic_vector(to_unsigned( 97,8)),
			12305 => std_logic_vector(to_unsigned( 160,8)),
			12306 => std_logic_vector(to_unsigned( 64,8)),
			12307 => std_logic_vector(to_unsigned( 112,8)),
			12308 => std_logic_vector(to_unsigned( 74,8)),
			12309 => std_logic_vector(to_unsigned( 254,8)),
			12310 => std_logic_vector(to_unsigned( 146,8)),
			12311 => std_logic_vector(to_unsigned( 4,8)),
			12312 => std_logic_vector(to_unsigned( 20,8)),
			12313 => std_logic_vector(to_unsigned( 248,8)),
			12314 => std_logic_vector(to_unsigned( 180,8)),
			12315 => std_logic_vector(to_unsigned( 174,8)),
			12316 => std_logic_vector(to_unsigned( 175,8)),
			12317 => std_logic_vector(to_unsigned( 37,8)),
			12318 => std_logic_vector(to_unsigned( 254,8)),
			12319 => std_logic_vector(to_unsigned( 253,8)),
			12320 => std_logic_vector(to_unsigned( 207,8)),
			12321 => std_logic_vector(to_unsigned( 217,8)),
			12322 => std_logic_vector(to_unsigned( 68,8)),
			12323 => std_logic_vector(to_unsigned( 126,8)),
			12324 => std_logic_vector(to_unsigned( 247,8)),
			12325 => std_logic_vector(to_unsigned( 130,8)),
			12326 => std_logic_vector(to_unsigned( 200,8)),
			12327 => std_logic_vector(to_unsigned( 128,8)),
			12328 => std_logic_vector(to_unsigned( 110,8)),
			12329 => std_logic_vector(to_unsigned( 42,8)),
			12330 => std_logic_vector(to_unsigned( 231,8)),
			12331 => std_logic_vector(to_unsigned( 168,8)),
			12332 => std_logic_vector(to_unsigned( 212,8)),
			12333 => std_logic_vector(to_unsigned( 104,8)),
			12334 => std_logic_vector(to_unsigned( 189,8)),
			12335 => std_logic_vector(to_unsigned( 58,8)),
			12336 => std_logic_vector(to_unsigned( 110,8)),
			12337 => std_logic_vector(to_unsigned( 250,8)),
			12338 => std_logic_vector(to_unsigned( 156,8)),
			12339 => std_logic_vector(to_unsigned( 92,8)),
			12340 => std_logic_vector(to_unsigned( 168,8)),
			12341 => std_logic_vector(to_unsigned( 215,8)),
			12342 => std_logic_vector(to_unsigned( 217,8)),
			12343 => std_logic_vector(to_unsigned( 76,8)),
			12344 => std_logic_vector(to_unsigned( 58,8)),
			12345 => std_logic_vector(to_unsigned( 131,8)),
			12346 => std_logic_vector(to_unsigned( 125,8)),
			12347 => std_logic_vector(to_unsigned( 0,8)),
			12348 => std_logic_vector(to_unsigned( 37,8)),
			12349 => std_logic_vector(to_unsigned( 169,8)),
			12350 => std_logic_vector(to_unsigned( 145,8)),
			12351 => std_logic_vector(to_unsigned( 75,8)),
			12352 => std_logic_vector(to_unsigned( 155,8)),
			12353 => std_logic_vector(to_unsigned( 65,8)),
			12354 => std_logic_vector(to_unsigned( 101,8)),
			12355 => std_logic_vector(to_unsigned( 212,8)),
			12356 => std_logic_vector(to_unsigned( 224,8)),
			12357 => std_logic_vector(to_unsigned( 193,8)),
			12358 => std_logic_vector(to_unsigned( 53,8)),
			12359 => std_logic_vector(to_unsigned( 249,8)),
			12360 => std_logic_vector(to_unsigned( 121,8)),
			12361 => std_logic_vector(to_unsigned( 115,8)),
			12362 => std_logic_vector(to_unsigned( 37,8)),
			12363 => std_logic_vector(to_unsigned( 255,8)),
			12364 => std_logic_vector(to_unsigned( 234,8)),
			12365 => std_logic_vector(to_unsigned( 232,8)),
			12366 => std_logic_vector(to_unsigned( 31,8)),
			12367 => std_logic_vector(to_unsigned( 81,8)),
			12368 => std_logic_vector(to_unsigned( 190,8)),
			12369 => std_logic_vector(to_unsigned( 69,8)),
			12370 => std_logic_vector(to_unsigned( 80,8)),
			12371 => std_logic_vector(to_unsigned( 31,8)),
			12372 => std_logic_vector(to_unsigned( 213,8)),
			12373 => std_logic_vector(to_unsigned( 130,8)),
			12374 => std_logic_vector(to_unsigned( 212,8)),
			12375 => std_logic_vector(to_unsigned( 16,8)),
			12376 => std_logic_vector(to_unsigned( 5,8)),
			12377 => std_logic_vector(to_unsigned( 168,8)),
			12378 => std_logic_vector(to_unsigned( 59,8)),
			12379 => std_logic_vector(to_unsigned( 56,8)),
			12380 => std_logic_vector(to_unsigned( 3,8)),
			12381 => std_logic_vector(to_unsigned( 35,8)),
			12382 => std_logic_vector(to_unsigned( 205,8)),
			12383 => std_logic_vector(to_unsigned( 180,8)),
			12384 => std_logic_vector(to_unsigned( 121,8)),
			12385 => std_logic_vector(to_unsigned( 169,8)),
			12386 => std_logic_vector(to_unsigned( 218,8)),
			12387 => std_logic_vector(to_unsigned( 27,8)),
			12388 => std_logic_vector(to_unsigned( 212,8)),
			12389 => std_logic_vector(to_unsigned( 157,8)),
			12390 => std_logic_vector(to_unsigned( 245,8)),
			12391 => std_logic_vector(to_unsigned( 59,8)),
			12392 => std_logic_vector(to_unsigned( 240,8)),
			12393 => std_logic_vector(to_unsigned( 174,8)),
			12394 => std_logic_vector(to_unsigned( 229,8)),
			12395 => std_logic_vector(to_unsigned( 151,8)),
			12396 => std_logic_vector(to_unsigned( 42,8)),
			12397 => std_logic_vector(to_unsigned( 101,8)),
			12398 => std_logic_vector(to_unsigned( 29,8)),
			12399 => std_logic_vector(to_unsigned( 252,8)),
			12400 => std_logic_vector(to_unsigned( 183,8)),
			12401 => std_logic_vector(to_unsigned( 71,8)),
			12402 => std_logic_vector(to_unsigned( 235,8)),
			12403 => std_logic_vector(to_unsigned( 172,8)),
			12404 => std_logic_vector(to_unsigned( 34,8)),
			12405 => std_logic_vector(to_unsigned( 63,8)),
			12406 => std_logic_vector(to_unsigned( 3,8)),
			12407 => std_logic_vector(to_unsigned( 26,8)),
			12408 => std_logic_vector(to_unsigned( 125,8)),
			12409 => std_logic_vector(to_unsigned( 51,8)),
			12410 => std_logic_vector(to_unsigned( 202,8)),
			12411 => std_logic_vector(to_unsigned( 8,8)),
			12412 => std_logic_vector(to_unsigned( 118,8)),
			12413 => std_logic_vector(to_unsigned( 148,8)),
			12414 => std_logic_vector(to_unsigned( 147,8)),
			12415 => std_logic_vector(to_unsigned( 199,8)),
			12416 => std_logic_vector(to_unsigned( 243,8)),
			12417 => std_logic_vector(to_unsigned( 13,8)),
			12418 => std_logic_vector(to_unsigned( 222,8)),
			12419 => std_logic_vector(to_unsigned( 64,8)),
			12420 => std_logic_vector(to_unsigned( 222,8)),
			12421 => std_logic_vector(to_unsigned( 214,8)),
			12422 => std_logic_vector(to_unsigned( 39,8)),
			12423 => std_logic_vector(to_unsigned( 219,8)),
			12424 => std_logic_vector(to_unsigned( 57,8)),
			12425 => std_logic_vector(to_unsigned( 136,8)),
			12426 => std_logic_vector(to_unsigned( 106,8)),
			12427 => std_logic_vector(to_unsigned( 40,8)),
			12428 => std_logic_vector(to_unsigned( 28,8)),
			12429 => std_logic_vector(to_unsigned( 129,8)),
			12430 => std_logic_vector(to_unsigned( 191,8)),
			12431 => std_logic_vector(to_unsigned( 193,8)),
			12432 => std_logic_vector(to_unsigned( 69,8)),
			12433 => std_logic_vector(to_unsigned( 78,8)),
			12434 => std_logic_vector(to_unsigned( 55,8)),
			12435 => std_logic_vector(to_unsigned( 173,8)),
			12436 => std_logic_vector(to_unsigned( 1,8)),
			12437 => std_logic_vector(to_unsigned( 213,8)),
			12438 => std_logic_vector(to_unsigned( 247,8)),
			12439 => std_logic_vector(to_unsigned( 221,8)),
			12440 => std_logic_vector(to_unsigned( 189,8)),
			12441 => std_logic_vector(to_unsigned( 22,8)),
			12442 => std_logic_vector(to_unsigned( 234,8)),
			12443 => std_logic_vector(to_unsigned( 220,8)),
			12444 => std_logic_vector(to_unsigned( 93,8)),
			12445 => std_logic_vector(to_unsigned( 212,8)),
			12446 => std_logic_vector(to_unsigned( 192,8)),
			12447 => std_logic_vector(to_unsigned( 143,8)),
			12448 => std_logic_vector(to_unsigned( 167,8)),
			12449 => std_logic_vector(to_unsigned( 219,8)),
			12450 => std_logic_vector(to_unsigned( 205,8)),
			12451 => std_logic_vector(to_unsigned( 9,8)),
			12452 => std_logic_vector(to_unsigned( 92,8)),
			12453 => std_logic_vector(to_unsigned( 181,8)),
			12454 => std_logic_vector(to_unsigned( 54,8)),
			12455 => std_logic_vector(to_unsigned( 15,8)),
			12456 => std_logic_vector(to_unsigned( 142,8)),
			12457 => std_logic_vector(to_unsigned( 103,8)),
			12458 => std_logic_vector(to_unsigned( 187,8)),
			12459 => std_logic_vector(to_unsigned( 106,8)),
			12460 => std_logic_vector(to_unsigned( 246,8)),
			12461 => std_logic_vector(to_unsigned( 130,8)),
			12462 => std_logic_vector(to_unsigned( 91,8)),
			12463 => std_logic_vector(to_unsigned( 171,8)),
			12464 => std_logic_vector(to_unsigned( 98,8)),
			12465 => std_logic_vector(to_unsigned( 152,8)),
			12466 => std_logic_vector(to_unsigned( 61,8)),
			12467 => std_logic_vector(to_unsigned( 232,8)),
			12468 => std_logic_vector(to_unsigned( 225,8)),
			12469 => std_logic_vector(to_unsigned( 243,8)),
			12470 => std_logic_vector(to_unsigned( 121,8)),
			12471 => std_logic_vector(to_unsigned( 218,8)),
			12472 => std_logic_vector(to_unsigned( 118,8)),
			12473 => std_logic_vector(to_unsigned( 68,8)),
			12474 => std_logic_vector(to_unsigned( 209,8)),
			12475 => std_logic_vector(to_unsigned( 194,8)),
			12476 => std_logic_vector(to_unsigned( 93,8)),
			12477 => std_logic_vector(to_unsigned( 114,8)),
			12478 => std_logic_vector(to_unsigned( 242,8)),
			12479 => std_logic_vector(to_unsigned( 33,8)),
			12480 => std_logic_vector(to_unsigned( 250,8)),
			12481 => std_logic_vector(to_unsigned( 247,8)),
			12482 => std_logic_vector(to_unsigned( 71,8)),
			12483 => std_logic_vector(to_unsigned( 147,8)),
			12484 => std_logic_vector(to_unsigned( 86,8)),
			12485 => std_logic_vector(to_unsigned( 146,8)),
			12486 => std_logic_vector(to_unsigned( 66,8)),
			12487 => std_logic_vector(to_unsigned( 75,8)),
			12488 => std_logic_vector(to_unsigned( 160,8)),
			12489 => std_logic_vector(to_unsigned( 35,8)),
			12490 => std_logic_vector(to_unsigned( 212,8)),
			12491 => std_logic_vector(to_unsigned( 44,8)),
			12492 => std_logic_vector(to_unsigned( 183,8)),
			12493 => std_logic_vector(to_unsigned( 196,8)),
			12494 => std_logic_vector(to_unsigned( 188,8)),
			12495 => std_logic_vector(to_unsigned( 10,8)),
			12496 => std_logic_vector(to_unsigned( 233,8)),
			12497 => std_logic_vector(to_unsigned( 24,8)),
			12498 => std_logic_vector(to_unsigned( 2,8)),
			12499 => std_logic_vector(to_unsigned( 247,8)),
			12500 => std_logic_vector(to_unsigned( 150,8)),
			12501 => std_logic_vector(to_unsigned( 248,8)),
			12502 => std_logic_vector(to_unsigned( 231,8)),
			12503 => std_logic_vector(to_unsigned( 37,8)),
			12504 => std_logic_vector(to_unsigned( 189,8)),
			12505 => std_logic_vector(to_unsigned( 120,8)),
			12506 => std_logic_vector(to_unsigned( 99,8)),
			12507 => std_logic_vector(to_unsigned( 152,8)),
			12508 => std_logic_vector(to_unsigned( 247,8)),
			12509 => std_logic_vector(to_unsigned( 226,8)),
			12510 => std_logic_vector(to_unsigned( 80,8)),
			12511 => std_logic_vector(to_unsigned( 193,8)),
			12512 => std_logic_vector(to_unsigned( 248,8)),
			12513 => std_logic_vector(to_unsigned( 89,8)),
			12514 => std_logic_vector(to_unsigned( 119,8)),
			12515 => std_logic_vector(to_unsigned( 172,8)),
			12516 => std_logic_vector(to_unsigned( 143,8)),
			12517 => std_logic_vector(to_unsigned( 244,8)),
			12518 => std_logic_vector(to_unsigned( 39,8)),
			12519 => std_logic_vector(to_unsigned( 99,8)),
			12520 => std_logic_vector(to_unsigned( 52,8)),
			12521 => std_logic_vector(to_unsigned( 9,8)),
			12522 => std_logic_vector(to_unsigned( 246,8)),
			12523 => std_logic_vector(to_unsigned( 206,8)),
			12524 => std_logic_vector(to_unsigned( 67,8)),
			12525 => std_logic_vector(to_unsigned( 55,8)),
			12526 => std_logic_vector(to_unsigned( 81,8)),
			12527 => std_logic_vector(to_unsigned( 196,8)),
			12528 => std_logic_vector(to_unsigned( 223,8)),
			12529 => std_logic_vector(to_unsigned( 155,8)),
			12530 => std_logic_vector(to_unsigned( 116,8)),
			12531 => std_logic_vector(to_unsigned( 180,8)),
			12532 => std_logic_vector(to_unsigned( 66,8)),
			12533 => std_logic_vector(to_unsigned( 184,8)),
			12534 => std_logic_vector(to_unsigned( 238,8)),
			12535 => std_logic_vector(to_unsigned( 29,8)),
			12536 => std_logic_vector(to_unsigned( 232,8)),
			12537 => std_logic_vector(to_unsigned( 110,8)),
			12538 => std_logic_vector(to_unsigned( 200,8)),
			12539 => std_logic_vector(to_unsigned( 148,8)),
			12540 => std_logic_vector(to_unsigned( 179,8)),
			12541 => std_logic_vector(to_unsigned( 227,8)),
			12542 => std_logic_vector(to_unsigned( 94,8)),
			12543 => std_logic_vector(to_unsigned( 66,8)),
			12544 => std_logic_vector(to_unsigned( 29,8)),
			12545 => std_logic_vector(to_unsigned( 120,8)),
			12546 => std_logic_vector(to_unsigned( 199,8)),
			12547 => std_logic_vector(to_unsigned( 122,8)),
			12548 => std_logic_vector(to_unsigned( 85,8)),
			12549 => std_logic_vector(to_unsigned( 186,8)),
			12550 => std_logic_vector(to_unsigned( 244,8)),
			12551 => std_logic_vector(to_unsigned( 72,8)),
			12552 => std_logic_vector(to_unsigned( 54,8)),
			12553 => std_logic_vector(to_unsigned( 182,8)),
			12554 => std_logic_vector(to_unsigned( 225,8)),
			12555 => std_logic_vector(to_unsigned( 226,8)),
			12556 => std_logic_vector(to_unsigned( 165,8)),
			12557 => std_logic_vector(to_unsigned( 132,8)),
			12558 => std_logic_vector(to_unsigned( 96,8)),
			12559 => std_logic_vector(to_unsigned( 43,8)),
			12560 => std_logic_vector(to_unsigned( 205,8)),
			12561 => std_logic_vector(to_unsigned( 206,8)),
			12562 => std_logic_vector(to_unsigned( 125,8)),
			12563 => std_logic_vector(to_unsigned( 70,8)),
			12564 => std_logic_vector(to_unsigned( 163,8)),
			12565 => std_logic_vector(to_unsigned( 67,8)),
			12566 => std_logic_vector(to_unsigned( 223,8)),
			12567 => std_logic_vector(to_unsigned( 173,8)),
			12568 => std_logic_vector(to_unsigned( 188,8)),
			12569 => std_logic_vector(to_unsigned( 2,8)),
			12570 => std_logic_vector(to_unsigned( 29,8)),
			12571 => std_logic_vector(to_unsigned( 43,8)),
			12572 => std_logic_vector(to_unsigned( 107,8)),
			12573 => std_logic_vector(to_unsigned( 105,8)),
			12574 => std_logic_vector(to_unsigned( 13,8)),
			12575 => std_logic_vector(to_unsigned( 60,8)),
			12576 => std_logic_vector(to_unsigned( 191,8)),
			12577 => std_logic_vector(to_unsigned( 23,8)),
			12578 => std_logic_vector(to_unsigned( 20,8)),
			12579 => std_logic_vector(to_unsigned( 157,8)),
			12580 => std_logic_vector(to_unsigned( 169,8)),
			12581 => std_logic_vector(to_unsigned( 207,8)),
			12582 => std_logic_vector(to_unsigned( 235,8)),
			12583 => std_logic_vector(to_unsigned( 220,8)),
			12584 => std_logic_vector(to_unsigned( 187,8)),
			12585 => std_logic_vector(to_unsigned( 183,8)),
			12586 => std_logic_vector(to_unsigned( 162,8)),
			12587 => std_logic_vector(to_unsigned( 20,8)),
			12588 => std_logic_vector(to_unsigned( 190,8)),
			12589 => std_logic_vector(to_unsigned( 179,8)),
			12590 => std_logic_vector(to_unsigned( 8,8)),
			12591 => std_logic_vector(to_unsigned( 222,8)),
			12592 => std_logic_vector(to_unsigned( 86,8)),
			12593 => std_logic_vector(to_unsigned( 199,8)),
			12594 => std_logic_vector(to_unsigned( 76,8)),
			12595 => std_logic_vector(to_unsigned( 242,8)),
			12596 => std_logic_vector(to_unsigned( 85,8)),
			12597 => std_logic_vector(to_unsigned( 166,8)),
			12598 => std_logic_vector(to_unsigned( 210,8)),
			12599 => std_logic_vector(to_unsigned( 213,8)),
			12600 => std_logic_vector(to_unsigned( 215,8)),
			12601 => std_logic_vector(to_unsigned( 110,8)),
			12602 => std_logic_vector(to_unsigned( 108,8)),
			12603 => std_logic_vector(to_unsigned( 169,8)),
			12604 => std_logic_vector(to_unsigned( 231,8)),
			12605 => std_logic_vector(to_unsigned( 98,8)),
			12606 => std_logic_vector(to_unsigned( 9,8)),
			12607 => std_logic_vector(to_unsigned( 253,8)),
			12608 => std_logic_vector(to_unsigned( 202,8)),
			12609 => std_logic_vector(to_unsigned( 153,8)),
			12610 => std_logic_vector(to_unsigned( 44,8)),
			12611 => std_logic_vector(to_unsigned( 154,8)),
			12612 => std_logic_vector(to_unsigned( 25,8)),
			12613 => std_logic_vector(to_unsigned( 82,8)),
			12614 => std_logic_vector(to_unsigned( 218,8)),
			12615 => std_logic_vector(to_unsigned( 93,8)),
			12616 => std_logic_vector(to_unsigned( 201,8)),
			12617 => std_logic_vector(to_unsigned( 252,8)),
			12618 => std_logic_vector(to_unsigned( 146,8)),
			12619 => std_logic_vector(to_unsigned( 238,8)),
			12620 => std_logic_vector(to_unsigned( 125,8)),
			12621 => std_logic_vector(to_unsigned( 46,8)),
			12622 => std_logic_vector(to_unsigned( 195,8)),
			12623 => std_logic_vector(to_unsigned( 168,8)),
			12624 => std_logic_vector(to_unsigned( 211,8)),
			12625 => std_logic_vector(to_unsigned( 111,8)),
			12626 => std_logic_vector(to_unsigned( 254,8)),
			12627 => std_logic_vector(to_unsigned( 224,8)),
			12628 => std_logic_vector(to_unsigned( 142,8)),
			12629 => std_logic_vector(to_unsigned( 15,8)),
			12630 => std_logic_vector(to_unsigned( 231,8)),
			12631 => std_logic_vector(to_unsigned( 62,8)),
			12632 => std_logic_vector(to_unsigned( 78,8)),
			12633 => std_logic_vector(to_unsigned( 104,8)),
			12634 => std_logic_vector(to_unsigned( 237,8)),
			12635 => std_logic_vector(to_unsigned( 135,8)),
			12636 => std_logic_vector(to_unsigned( 231,8)),
			12637 => std_logic_vector(to_unsigned( 85,8)),
			12638 => std_logic_vector(to_unsigned( 184,8)),
			12639 => std_logic_vector(to_unsigned( 14,8)),
			12640 => std_logic_vector(to_unsigned( 172,8)),
			12641 => std_logic_vector(to_unsigned( 105,8)),
			12642 => std_logic_vector(to_unsigned( 165,8)),
			12643 => std_logic_vector(to_unsigned( 243,8)),
			12644 => std_logic_vector(to_unsigned( 220,8)),
			12645 => std_logic_vector(to_unsigned( 32,8)),
			12646 => std_logic_vector(to_unsigned( 149,8)),
			12647 => std_logic_vector(to_unsigned( 194,8)),
			12648 => std_logic_vector(to_unsigned( 150,8)),
			12649 => std_logic_vector(to_unsigned( 47,8)),
			12650 => std_logic_vector(to_unsigned( 82,8)),
			12651 => std_logic_vector(to_unsigned( 81,8)),
			12652 => std_logic_vector(to_unsigned( 167,8)),
			12653 => std_logic_vector(to_unsigned( 76,8)),
			12654 => std_logic_vector(to_unsigned( 208,8)),
			12655 => std_logic_vector(to_unsigned( 228,8)),
			12656 => std_logic_vector(to_unsigned( 235,8)),
			12657 => std_logic_vector(to_unsigned( 237,8)),
			12658 => std_logic_vector(to_unsigned( 233,8)),
			12659 => std_logic_vector(to_unsigned( 223,8)),
			12660 => std_logic_vector(to_unsigned( 226,8)),
			12661 => std_logic_vector(to_unsigned( 144,8)),
			12662 => std_logic_vector(to_unsigned( 126,8)),
			12663 => std_logic_vector(to_unsigned( 86,8)),
			12664 => std_logic_vector(to_unsigned( 142,8)),
			12665 => std_logic_vector(to_unsigned( 165,8)),
			12666 => std_logic_vector(to_unsigned( 117,8)),
			12667 => std_logic_vector(to_unsigned( 142,8)),
			12668 => std_logic_vector(to_unsigned( 145,8)),
			12669 => std_logic_vector(to_unsigned( 229,8)),
			12670 => std_logic_vector(to_unsigned( 81,8)),
			12671 => std_logic_vector(to_unsigned( 186,8)),
			12672 => std_logic_vector(to_unsigned( 136,8)),
			12673 => std_logic_vector(to_unsigned( 194,8)),
			12674 => std_logic_vector(to_unsigned( 56,8)),
			12675 => std_logic_vector(to_unsigned( 83,8)),
			12676 => std_logic_vector(to_unsigned( 156,8)),
			12677 => std_logic_vector(to_unsigned( 219,8)),
			12678 => std_logic_vector(to_unsigned( 99,8)),
			12679 => std_logic_vector(to_unsigned( 80,8)),
			12680 => std_logic_vector(to_unsigned( 114,8)),
			12681 => std_logic_vector(to_unsigned( 97,8)),
			12682 => std_logic_vector(to_unsigned( 252,8)),
			12683 => std_logic_vector(to_unsigned( 186,8)),
			12684 => std_logic_vector(to_unsigned( 254,8)),
			12685 => std_logic_vector(to_unsigned( 19,8)),
			12686 => std_logic_vector(to_unsigned( 15,8)),
			12687 => std_logic_vector(to_unsigned( 252,8)),
			12688 => std_logic_vector(to_unsigned( 29,8)),
			12689 => std_logic_vector(to_unsigned( 64,8)),
			12690 => std_logic_vector(to_unsigned( 104,8)),
			12691 => std_logic_vector(to_unsigned( 22,8)),
			12692 => std_logic_vector(to_unsigned( 156,8)),
			12693 => std_logic_vector(to_unsigned( 155,8)),
			12694 => std_logic_vector(to_unsigned( 212,8)),
			12695 => std_logic_vector(to_unsigned( 42,8)),
			12696 => std_logic_vector(to_unsigned( 40,8)),
			12697 => std_logic_vector(to_unsigned( 165,8)),
			12698 => std_logic_vector(to_unsigned( 69,8)),
			12699 => std_logic_vector(to_unsigned( 177,8)),
			12700 => std_logic_vector(to_unsigned( 1,8)),
			12701 => std_logic_vector(to_unsigned( 170,8)),
			12702 => std_logic_vector(to_unsigned( 227,8)),
			12703 => std_logic_vector(to_unsigned( 184,8)),
			12704 => std_logic_vector(to_unsigned( 63,8)),
			12705 => std_logic_vector(to_unsigned( 46,8)),
			12706 => std_logic_vector(to_unsigned( 149,8)),
			12707 => std_logic_vector(to_unsigned( 0,8)),
			12708 => std_logic_vector(to_unsigned( 225,8)),
			12709 => std_logic_vector(to_unsigned( 63,8)),
			12710 => std_logic_vector(to_unsigned( 100,8)),
			12711 => std_logic_vector(to_unsigned( 14,8)),
			12712 => std_logic_vector(to_unsigned( 35,8)),
			12713 => std_logic_vector(to_unsigned( 235,8)),
			12714 => std_logic_vector(to_unsigned( 27,8)),
			12715 => std_logic_vector(to_unsigned( 137,8)),
			12716 => std_logic_vector(to_unsigned( 240,8)),
			12717 => std_logic_vector(to_unsigned( 145,8)),
			12718 => std_logic_vector(to_unsigned( 171,8)),
			12719 => std_logic_vector(to_unsigned( 117,8)),
			12720 => std_logic_vector(to_unsigned( 188,8)),
			12721 => std_logic_vector(to_unsigned( 229,8)),
			12722 => std_logic_vector(to_unsigned( 234,8)),
			12723 => std_logic_vector(to_unsigned( 96,8)),
			12724 => std_logic_vector(to_unsigned( 80,8)),
			12725 => std_logic_vector(to_unsigned( 18,8)),
			12726 => std_logic_vector(to_unsigned( 107,8)),
			12727 => std_logic_vector(to_unsigned( 28,8)),
			12728 => std_logic_vector(to_unsigned( 7,8)),
			12729 => std_logic_vector(to_unsigned( 0,8)),
			12730 => std_logic_vector(to_unsigned( 9,8)),
			12731 => std_logic_vector(to_unsigned( 143,8)),
			12732 => std_logic_vector(to_unsigned( 76,8)),
			12733 => std_logic_vector(to_unsigned( 203,8)),
			12734 => std_logic_vector(to_unsigned( 26,8)),
			12735 => std_logic_vector(to_unsigned( 184,8)),
			12736 => std_logic_vector(to_unsigned( 200,8)),
			12737 => std_logic_vector(to_unsigned( 186,8)),
			12738 => std_logic_vector(to_unsigned( 31,8)),
			12739 => std_logic_vector(to_unsigned( 114,8)),
			12740 => std_logic_vector(to_unsigned( 54,8)),
			12741 => std_logic_vector(to_unsigned( 132,8)),
			12742 => std_logic_vector(to_unsigned( 101,8)),
			12743 => std_logic_vector(to_unsigned( 146,8)),
			12744 => std_logic_vector(to_unsigned( 211,8)),
			12745 => std_logic_vector(to_unsigned( 225,8)),
			12746 => std_logic_vector(to_unsigned( 191,8)),
			12747 => std_logic_vector(to_unsigned( 175,8)),
			12748 => std_logic_vector(to_unsigned( 63,8)),
			12749 => std_logic_vector(to_unsigned( 222,8)),
			12750 => std_logic_vector(to_unsigned( 49,8)),
			12751 => std_logic_vector(to_unsigned( 15,8)),
			12752 => std_logic_vector(to_unsigned( 79,8)),
			12753 => std_logic_vector(to_unsigned( 104,8)),
			12754 => std_logic_vector(to_unsigned( 97,8)),
			12755 => std_logic_vector(to_unsigned( 7,8)),
			12756 => std_logic_vector(to_unsigned( 89,8)),
			12757 => std_logic_vector(to_unsigned( 120,8)),
			12758 => std_logic_vector(to_unsigned( 172,8)),
			12759 => std_logic_vector(to_unsigned( 39,8)),
			12760 => std_logic_vector(to_unsigned( 132,8)),
			12761 => std_logic_vector(to_unsigned( 100,8)),
			12762 => std_logic_vector(to_unsigned( 160,8)),
			12763 => std_logic_vector(to_unsigned( 3,8)),
			12764 => std_logic_vector(to_unsigned( 220,8)),
			12765 => std_logic_vector(to_unsigned( 75,8)),
			12766 => std_logic_vector(to_unsigned( 247,8)),
			12767 => std_logic_vector(to_unsigned( 122,8)),
			12768 => std_logic_vector(to_unsigned( 197,8)),
			12769 => std_logic_vector(to_unsigned( 10,8)),
			12770 => std_logic_vector(to_unsigned( 110,8)),
			12771 => std_logic_vector(to_unsigned( 40,8)),
			12772 => std_logic_vector(to_unsigned( 76,8)),
			12773 => std_logic_vector(to_unsigned( 149,8)),
			12774 => std_logic_vector(to_unsigned( 209,8)),
			12775 => std_logic_vector(to_unsigned( 90,8)),
			12776 => std_logic_vector(to_unsigned( 231,8)),
			12777 => std_logic_vector(to_unsigned( 202,8)),
			12778 => std_logic_vector(to_unsigned( 176,8)),
			12779 => std_logic_vector(to_unsigned( 254,8)),
			12780 => std_logic_vector(to_unsigned( 122,8)),
			12781 => std_logic_vector(to_unsigned( 43,8)),
			12782 => std_logic_vector(to_unsigned( 94,8)),
			12783 => std_logic_vector(to_unsigned( 157,8)),
			12784 => std_logic_vector(to_unsigned( 54,8)),
			12785 => std_logic_vector(to_unsigned( 123,8)),
			12786 => std_logic_vector(to_unsigned( 230,8)),
			12787 => std_logic_vector(to_unsigned( 242,8)),
			12788 => std_logic_vector(to_unsigned( 168,8)),
			12789 => std_logic_vector(to_unsigned( 65,8)),
			12790 => std_logic_vector(to_unsigned( 145,8)),
			12791 => std_logic_vector(to_unsigned( 229,8)),
			12792 => std_logic_vector(to_unsigned( 33,8)),
			12793 => std_logic_vector(to_unsigned( 182,8)),
			12794 => std_logic_vector(to_unsigned( 12,8)),
			12795 => std_logic_vector(to_unsigned( 133,8)),
			12796 => std_logic_vector(to_unsigned( 0,8)),
			12797 => std_logic_vector(to_unsigned( 134,8)),
			12798 => std_logic_vector(to_unsigned( 108,8)),
			12799 => std_logic_vector(to_unsigned( 167,8)),
			12800 => std_logic_vector(to_unsigned( 197,8)),
			12801 => std_logic_vector(to_unsigned( 135,8)),
			12802 => std_logic_vector(to_unsigned( 214,8)),
			12803 => std_logic_vector(to_unsigned( 242,8)),
			12804 => std_logic_vector(to_unsigned( 115,8)),
			12805 => std_logic_vector(to_unsigned( 172,8)),
			12806 => std_logic_vector(to_unsigned( 20,8)),
			12807 => std_logic_vector(to_unsigned( 58,8)),
			12808 => std_logic_vector(to_unsigned( 140,8)),
			12809 => std_logic_vector(to_unsigned( 84,8)),
			12810 => std_logic_vector(to_unsigned( 200,8)),
			12811 => std_logic_vector(to_unsigned( 85,8)),
			12812 => std_logic_vector(to_unsigned( 154,8)),
			12813 => std_logic_vector(to_unsigned( 34,8)),
			12814 => std_logic_vector(to_unsigned( 181,8)),
			12815 => std_logic_vector(to_unsigned( 128,8)),
			12816 => std_logic_vector(to_unsigned( 78,8)),
			12817 => std_logic_vector(to_unsigned( 235,8)),
			12818 => std_logic_vector(to_unsigned( 80,8)),
			12819 => std_logic_vector(to_unsigned( 72,8)),
			12820 => std_logic_vector(to_unsigned( 28,8)),
			12821 => std_logic_vector(to_unsigned( 221,8)),
			12822 => std_logic_vector(to_unsigned( 250,8)),
			12823 => std_logic_vector(to_unsigned( 148,8)),
			12824 => std_logic_vector(to_unsigned( 10,8)),
			12825 => std_logic_vector(to_unsigned( 240,8)),
			12826 => std_logic_vector(to_unsigned( 236,8)),
			12827 => std_logic_vector(to_unsigned( 231,8)),
			12828 => std_logic_vector(to_unsigned( 183,8)),
			12829 => std_logic_vector(to_unsigned( 166,8)),
			12830 => std_logic_vector(to_unsigned( 65,8)),
			12831 => std_logic_vector(to_unsigned( 253,8)),
			12832 => std_logic_vector(to_unsigned( 128,8)),
			12833 => std_logic_vector(to_unsigned( 212,8)),
			12834 => std_logic_vector(to_unsigned( 101,8)),
			12835 => std_logic_vector(to_unsigned( 14,8)),
			12836 => std_logic_vector(to_unsigned( 72,8)),
			12837 => std_logic_vector(to_unsigned( 1,8)),
			12838 => std_logic_vector(to_unsigned( 45,8)),
			12839 => std_logic_vector(to_unsigned( 13,8)),
			12840 => std_logic_vector(to_unsigned( 178,8)),
			12841 => std_logic_vector(to_unsigned( 56,8)),
			12842 => std_logic_vector(to_unsigned( 153,8)),
			12843 => std_logic_vector(to_unsigned( 9,8)),
			12844 => std_logic_vector(to_unsigned( 224,8)),
			12845 => std_logic_vector(to_unsigned( 15,8)),
			12846 => std_logic_vector(to_unsigned( 45,8)),
			12847 => std_logic_vector(to_unsigned( 78,8)),
			12848 => std_logic_vector(to_unsigned( 187,8)),
			12849 => std_logic_vector(to_unsigned( 225,8)),
			12850 => std_logic_vector(to_unsigned( 243,8)),
			12851 => std_logic_vector(to_unsigned( 157,8)),
			12852 => std_logic_vector(to_unsigned( 192,8)),
			12853 => std_logic_vector(to_unsigned( 79,8)),
			12854 => std_logic_vector(to_unsigned( 81,8)),
			12855 => std_logic_vector(to_unsigned( 18,8)),
			12856 => std_logic_vector(to_unsigned( 233,8)),
			12857 => std_logic_vector(to_unsigned( 252,8)),
			12858 => std_logic_vector(to_unsigned( 171,8)),
			12859 => std_logic_vector(to_unsigned( 64,8)),
			12860 => std_logic_vector(to_unsigned( 168,8)),
			12861 => std_logic_vector(to_unsigned( 228,8)),
			12862 => std_logic_vector(to_unsigned( 196,8)),
			12863 => std_logic_vector(to_unsigned( 147,8)),
			12864 => std_logic_vector(to_unsigned( 69,8)),
			12865 => std_logic_vector(to_unsigned( 71,8)),
			12866 => std_logic_vector(to_unsigned( 105,8)),
			12867 => std_logic_vector(to_unsigned( 200,8)),
			12868 => std_logic_vector(to_unsigned( 158,8)),
			12869 => std_logic_vector(to_unsigned( 177,8)),
			12870 => std_logic_vector(to_unsigned( 154,8)),
			12871 => std_logic_vector(to_unsigned( 167,8)),
			12872 => std_logic_vector(to_unsigned( 195,8)),
			12873 => std_logic_vector(to_unsigned( 94,8)),
			12874 => std_logic_vector(to_unsigned( 155,8)),
			12875 => std_logic_vector(to_unsigned( 94,8)),
			12876 => std_logic_vector(to_unsigned( 8,8)),
			12877 => std_logic_vector(to_unsigned( 222,8)),
			12878 => std_logic_vector(to_unsigned( 150,8)),
			12879 => std_logic_vector(to_unsigned( 32,8)),
			12880 => std_logic_vector(to_unsigned( 78,8)),
			12881 => std_logic_vector(to_unsigned( 238,8)),
			12882 => std_logic_vector(to_unsigned( 75,8)),
			12883 => std_logic_vector(to_unsigned( 83,8)),
			12884 => std_logic_vector(to_unsigned( 103,8)),
			12885 => std_logic_vector(to_unsigned( 109,8)),
			12886 => std_logic_vector(to_unsigned( 247,8)),
			12887 => std_logic_vector(to_unsigned( 235,8)),
			12888 => std_logic_vector(to_unsigned( 181,8)),
			12889 => std_logic_vector(to_unsigned( 2,8)),
			12890 => std_logic_vector(to_unsigned( 217,8)),
			12891 => std_logic_vector(to_unsigned( 242,8)),
			12892 => std_logic_vector(to_unsigned( 242,8)),
			12893 => std_logic_vector(to_unsigned( 35,8)),
			12894 => std_logic_vector(to_unsigned( 30,8)),
			12895 => std_logic_vector(to_unsigned( 18,8)),
			12896 => std_logic_vector(to_unsigned( 129,8)),
			12897 => std_logic_vector(to_unsigned( 235,8)),
			12898 => std_logic_vector(to_unsigned( 223,8)),
			12899 => std_logic_vector(to_unsigned( 69,8)),
			12900 => std_logic_vector(to_unsigned( 23,8)),
			12901 => std_logic_vector(to_unsigned( 171,8)),
			12902 => std_logic_vector(to_unsigned( 196,8)),
			12903 => std_logic_vector(to_unsigned( 129,8)),
			12904 => std_logic_vector(to_unsigned( 215,8)),
			12905 => std_logic_vector(to_unsigned( 50,8)),
			12906 => std_logic_vector(to_unsigned( 115,8)),
			12907 => std_logic_vector(to_unsigned( 228,8)),
			12908 => std_logic_vector(to_unsigned( 18,8)),
			12909 => std_logic_vector(to_unsigned( 171,8)),
			12910 => std_logic_vector(to_unsigned( 105,8)),
			12911 => std_logic_vector(to_unsigned( 64,8)),
			12912 => std_logic_vector(to_unsigned( 123,8)),
			12913 => std_logic_vector(to_unsigned( 98,8)),
			12914 => std_logic_vector(to_unsigned( 250,8)),
			12915 => std_logic_vector(to_unsigned( 25,8)),
			12916 => std_logic_vector(to_unsigned( 38,8)),
			12917 => std_logic_vector(to_unsigned( 178,8)),
			12918 => std_logic_vector(to_unsigned( 208,8)),
			12919 => std_logic_vector(to_unsigned( 88,8)),
			12920 => std_logic_vector(to_unsigned( 118,8)),
			12921 => std_logic_vector(to_unsigned( 12,8)),
			12922 => std_logic_vector(to_unsigned( 4,8)),
			12923 => std_logic_vector(to_unsigned( 253,8)),
			12924 => std_logic_vector(to_unsigned( 39,8)),
			12925 => std_logic_vector(to_unsigned( 48,8)),
			12926 => std_logic_vector(to_unsigned( 230,8)),
			12927 => std_logic_vector(to_unsigned( 194,8)),
			12928 => std_logic_vector(to_unsigned( 172,8)),
			12929 => std_logic_vector(to_unsigned( 40,8)),
			12930 => std_logic_vector(to_unsigned( 94,8)),
			12931 => std_logic_vector(to_unsigned( 102,8)),
			12932 => std_logic_vector(to_unsigned( 114,8)),
			12933 => std_logic_vector(to_unsigned( 139,8)),
			12934 => std_logic_vector(to_unsigned( 41,8)),
			12935 => std_logic_vector(to_unsigned( 163,8)),
			12936 => std_logic_vector(to_unsigned( 169,8)),
			12937 => std_logic_vector(to_unsigned( 195,8)),
			12938 => std_logic_vector(to_unsigned( 126,8)),
			12939 => std_logic_vector(to_unsigned( 6,8)),
			12940 => std_logic_vector(to_unsigned( 86,8)),
			12941 => std_logic_vector(to_unsigned( 173,8)),
			12942 => std_logic_vector(to_unsigned( 33,8)),
			12943 => std_logic_vector(to_unsigned( 226,8)),
			12944 => std_logic_vector(to_unsigned( 78,8)),
			12945 => std_logic_vector(to_unsigned( 90,8)),
			12946 => std_logic_vector(to_unsigned( 188,8)),
			12947 => std_logic_vector(to_unsigned( 168,8)),
			12948 => std_logic_vector(to_unsigned( 224,8)),
			12949 => std_logic_vector(to_unsigned( 181,8)),
			12950 => std_logic_vector(to_unsigned( 228,8)),
			12951 => std_logic_vector(to_unsigned( 141,8)),
			12952 => std_logic_vector(to_unsigned( 248,8)),
			12953 => std_logic_vector(to_unsigned( 24,8)),
			12954 => std_logic_vector(to_unsigned( 62,8)),
			12955 => std_logic_vector(to_unsigned( 173,8)),
			12956 => std_logic_vector(to_unsigned( 180,8)),
			12957 => std_logic_vector(to_unsigned( 61,8)),
			12958 => std_logic_vector(to_unsigned( 232,8)),
			12959 => std_logic_vector(to_unsigned( 1,8)),
			12960 => std_logic_vector(to_unsigned( 197,8)),
			12961 => std_logic_vector(to_unsigned( 107,8)),
			12962 => std_logic_vector(to_unsigned( 62,8)),
			12963 => std_logic_vector(to_unsigned( 198,8)),
			12964 => std_logic_vector(to_unsigned( 169,8)),
			12965 => std_logic_vector(to_unsigned( 86,8)),
			12966 => std_logic_vector(to_unsigned( 39,8)),
			12967 => std_logic_vector(to_unsigned( 8,8)),
			12968 => std_logic_vector(to_unsigned( 105,8)),
			12969 => std_logic_vector(to_unsigned( 111,8)),
			12970 => std_logic_vector(to_unsigned( 127,8)),
			12971 => std_logic_vector(to_unsigned( 41,8)),
			12972 => std_logic_vector(to_unsigned( 13,8)),
			12973 => std_logic_vector(to_unsigned( 49,8)),
			12974 => std_logic_vector(to_unsigned( 89,8)),
			12975 => std_logic_vector(to_unsigned( 22,8)),
			12976 => std_logic_vector(to_unsigned( 59,8)),
			12977 => std_logic_vector(to_unsigned( 99,8)),
			12978 => std_logic_vector(to_unsigned( 25,8)),
			12979 => std_logic_vector(to_unsigned( 184,8)),
			12980 => std_logic_vector(to_unsigned( 48,8)),
			12981 => std_logic_vector(to_unsigned( 218,8)),
			12982 => std_logic_vector(to_unsigned( 80,8)),
			12983 => std_logic_vector(to_unsigned( 65,8)),
			12984 => std_logic_vector(to_unsigned( 160,8)),
			12985 => std_logic_vector(to_unsigned( 75,8)),
			12986 => std_logic_vector(to_unsigned( 172,8)),
			12987 => std_logic_vector(to_unsigned( 250,8)),
			12988 => std_logic_vector(to_unsigned( 229,8)),
			12989 => std_logic_vector(to_unsigned( 76,8)),
			12990 => std_logic_vector(to_unsigned( 138,8)),
			12991 => std_logic_vector(to_unsigned( 223,8)),
			12992 => std_logic_vector(to_unsigned( 218,8)),
			12993 => std_logic_vector(to_unsigned( 83,8)),
			12994 => std_logic_vector(to_unsigned( 199,8)),
			12995 => std_logic_vector(to_unsigned( 211,8)),
			12996 => std_logic_vector(to_unsigned( 36,8)),
			12997 => std_logic_vector(to_unsigned( 202,8)),
			12998 => std_logic_vector(to_unsigned( 40,8)),
			12999 => std_logic_vector(to_unsigned( 48,8)),
			13000 => std_logic_vector(to_unsigned( 152,8)),
			13001 => std_logic_vector(to_unsigned( 3,8)),
			13002 => std_logic_vector(to_unsigned( 154,8)),
			13003 => std_logic_vector(to_unsigned( 171,8)),
			13004 => std_logic_vector(to_unsigned( 76,8)),
			13005 => std_logic_vector(to_unsigned( 161,8)),
			13006 => std_logic_vector(to_unsigned( 163,8)),
			13007 => std_logic_vector(to_unsigned( 227,8)),
			13008 => std_logic_vector(to_unsigned( 245,8)),
			13009 => std_logic_vector(to_unsigned( 214,8)),
			13010 => std_logic_vector(to_unsigned( 214,8)),
			13011 => std_logic_vector(to_unsigned( 110,8)),
			13012 => std_logic_vector(to_unsigned( 189,8)),
			13013 => std_logic_vector(to_unsigned( 208,8)),
			13014 => std_logic_vector(to_unsigned( 228,8)),
			13015 => std_logic_vector(to_unsigned( 208,8)),
			13016 => std_logic_vector(to_unsigned( 151,8)),
			13017 => std_logic_vector(to_unsigned( 78,8)),
			13018 => std_logic_vector(to_unsigned( 49,8)),
			13019 => std_logic_vector(to_unsigned( 5,8)),
			13020 => std_logic_vector(to_unsigned( 149,8)),
			13021 => std_logic_vector(to_unsigned( 239,8)),
			13022 => std_logic_vector(to_unsigned( 66,8)),
			13023 => std_logic_vector(to_unsigned( 253,8)),
			13024 => std_logic_vector(to_unsigned( 22,8)),
			13025 => std_logic_vector(to_unsigned( 200,8)),
			13026 => std_logic_vector(to_unsigned( 106,8)),
			13027 => std_logic_vector(to_unsigned( 84,8)),
			13028 => std_logic_vector(to_unsigned( 165,8)),
			13029 => std_logic_vector(to_unsigned( 129,8)),
			13030 => std_logic_vector(to_unsigned( 22,8)),
			13031 => std_logic_vector(to_unsigned( 77,8)),
			13032 => std_logic_vector(to_unsigned( 144,8)),
			13033 => std_logic_vector(to_unsigned( 218,8)),
			13034 => std_logic_vector(to_unsigned( 77,8)),
			13035 => std_logic_vector(to_unsigned( 153,8)),
			13036 => std_logic_vector(to_unsigned( 80,8)),
			13037 => std_logic_vector(to_unsigned( 245,8)),
			13038 => std_logic_vector(to_unsigned( 228,8)),
			13039 => std_logic_vector(to_unsigned( 9,8)),
			13040 => std_logic_vector(to_unsigned( 51,8)),
			13041 => std_logic_vector(to_unsigned( 124,8)),
			13042 => std_logic_vector(to_unsigned( 196,8)),
			13043 => std_logic_vector(to_unsigned( 154,8)),
			13044 => std_logic_vector(to_unsigned( 64,8)),
			13045 => std_logic_vector(to_unsigned( 194,8)),
			13046 => std_logic_vector(to_unsigned( 134,8)),
			13047 => std_logic_vector(to_unsigned( 234,8)),
			13048 => std_logic_vector(to_unsigned( 237,8)),
			13049 => std_logic_vector(to_unsigned( 99,8)),
			13050 => std_logic_vector(to_unsigned( 31,8)),
			13051 => std_logic_vector(to_unsigned( 137,8)),
			13052 => std_logic_vector(to_unsigned( 16,8)),
			13053 => std_logic_vector(to_unsigned( 89,8)),
			13054 => std_logic_vector(to_unsigned( 247,8)),
			13055 => std_logic_vector(to_unsigned( 88,8)),
			13056 => std_logic_vector(to_unsigned( 232,8)),
			13057 => std_logic_vector(to_unsigned( 57,8)),
			13058 => std_logic_vector(to_unsigned( 196,8)),
			13059 => std_logic_vector(to_unsigned( 134,8)),
			13060 => std_logic_vector(to_unsigned( 146,8)),
			13061 => std_logic_vector(to_unsigned( 96,8)),
			13062 => std_logic_vector(to_unsigned( 194,8)),
			13063 => std_logic_vector(to_unsigned( 185,8)),
			13064 => std_logic_vector(to_unsigned( 61,8)),
			13065 => std_logic_vector(to_unsigned( 23,8)),
			13066 => std_logic_vector(to_unsigned( 142,8)),
			13067 => std_logic_vector(to_unsigned( 131,8)),
			13068 => std_logic_vector(to_unsigned( 177,8)),
			13069 => std_logic_vector(to_unsigned( 221,8)),
			13070 => std_logic_vector(to_unsigned( 205,8)),
			13071 => std_logic_vector(to_unsigned( 5,8)),
			13072 => std_logic_vector(to_unsigned( 207,8)),
			13073 => std_logic_vector(to_unsigned( 253,8)),
			13074 => std_logic_vector(to_unsigned( 18,8)),
			13075 => std_logic_vector(to_unsigned( 28,8)),
			13076 => std_logic_vector(to_unsigned( 212,8)),
			13077 => std_logic_vector(to_unsigned( 93,8)),
			13078 => std_logic_vector(to_unsigned( 192,8)),
			13079 => std_logic_vector(to_unsigned( 29,8)),
			13080 => std_logic_vector(to_unsigned( 217,8)),
			13081 => std_logic_vector(to_unsigned( 175,8)),
			13082 => std_logic_vector(to_unsigned( 57,8)),
			13083 => std_logic_vector(to_unsigned( 184,8)),
			13084 => std_logic_vector(to_unsigned( 148,8)),
			13085 => std_logic_vector(to_unsigned( 17,8)),
			13086 => std_logic_vector(to_unsigned( 234,8)),
			13087 => std_logic_vector(to_unsigned( 133,8)),
			13088 => std_logic_vector(to_unsigned( 215,8)),
			13089 => std_logic_vector(to_unsigned( 15,8)),
			13090 => std_logic_vector(to_unsigned( 177,8)),
			13091 => std_logic_vector(to_unsigned( 234,8)),
			13092 => std_logic_vector(to_unsigned( 7,8)),
			13093 => std_logic_vector(to_unsigned( 155,8)),
			13094 => std_logic_vector(to_unsigned( 109,8)),
			13095 => std_logic_vector(to_unsigned( 155,8)),
			13096 => std_logic_vector(to_unsigned( 205,8)),
			13097 => std_logic_vector(to_unsigned( 86,8)),
			13098 => std_logic_vector(to_unsigned( 235,8)),
			13099 => std_logic_vector(to_unsigned( 170,8)),
			13100 => std_logic_vector(to_unsigned( 241,8)),
			13101 => std_logic_vector(to_unsigned( 250,8)),
			13102 => std_logic_vector(to_unsigned( 1,8)),
			13103 => std_logic_vector(to_unsigned( 41,8)),
			13104 => std_logic_vector(to_unsigned( 244,8)),
			13105 => std_logic_vector(to_unsigned( 142,8)),
			13106 => std_logic_vector(to_unsigned( 108,8)),
			13107 => std_logic_vector(to_unsigned( 165,8)),
			13108 => std_logic_vector(to_unsigned( 90,8)),
			13109 => std_logic_vector(to_unsigned( 239,8)),
			13110 => std_logic_vector(to_unsigned( 158,8)),
			13111 => std_logic_vector(to_unsigned( 22,8)),
			13112 => std_logic_vector(to_unsigned( 148,8)),
			13113 => std_logic_vector(to_unsigned( 174,8)),
			13114 => std_logic_vector(to_unsigned( 195,8)),
			13115 => std_logic_vector(to_unsigned( 45,8)),
			13116 => std_logic_vector(to_unsigned( 90,8)),
			13117 => std_logic_vector(to_unsigned( 157,8)),
			13118 => std_logic_vector(to_unsigned( 118,8)),
			13119 => std_logic_vector(to_unsigned( 181,8)),
			13120 => std_logic_vector(to_unsigned( 66,8)),
			13121 => std_logic_vector(to_unsigned( 245,8)),
			13122 => std_logic_vector(to_unsigned( 206,8)),
			13123 => std_logic_vector(to_unsigned( 80,8)),
			13124 => std_logic_vector(to_unsigned( 108,8)),
			13125 => std_logic_vector(to_unsigned( 83,8)),
			13126 => std_logic_vector(to_unsigned( 140,8)),
			13127 => std_logic_vector(to_unsigned( 196,8)),
			13128 => std_logic_vector(to_unsigned( 189,8)),
			13129 => std_logic_vector(to_unsigned( 149,8)),
			13130 => std_logic_vector(to_unsigned( 171,8)),
			13131 => std_logic_vector(to_unsigned( 86,8)),
			13132 => std_logic_vector(to_unsigned( 26,8)),
			13133 => std_logic_vector(to_unsigned( 64,8)),
			13134 => std_logic_vector(to_unsigned( 145,8)),
			13135 => std_logic_vector(to_unsigned( 126,8)),
			13136 => std_logic_vector(to_unsigned( 142,8)),
			13137 => std_logic_vector(to_unsigned( 180,8)),
			13138 => std_logic_vector(to_unsigned( 221,8)),
			13139 => std_logic_vector(to_unsigned( 216,8)),
			13140 => std_logic_vector(to_unsigned( 38,8)),
			13141 => std_logic_vector(to_unsigned( 222,8)),
			13142 => std_logic_vector(to_unsigned( 203,8)),
			13143 => std_logic_vector(to_unsigned( 156,8)),
			13144 => std_logic_vector(to_unsigned( 43,8)),
			13145 => std_logic_vector(to_unsigned( 32,8)),
			13146 => std_logic_vector(to_unsigned( 73,8)),
			13147 => std_logic_vector(to_unsigned( 155,8)),
			13148 => std_logic_vector(to_unsigned( 150,8)),
			13149 => std_logic_vector(to_unsigned( 249,8)),
			13150 => std_logic_vector(to_unsigned( 238,8)),
			13151 => std_logic_vector(to_unsigned( 42,8)),
			13152 => std_logic_vector(to_unsigned( 29,8)),
			13153 => std_logic_vector(to_unsigned( 119,8)),
			13154 => std_logic_vector(to_unsigned( 199,8)),
			13155 => std_logic_vector(to_unsigned( 133,8)),
			13156 => std_logic_vector(to_unsigned( 224,8)),
			13157 => std_logic_vector(to_unsigned( 40,8)),
			13158 => std_logic_vector(to_unsigned( 42,8)),
			13159 => std_logic_vector(to_unsigned( 191,8)),
			13160 => std_logic_vector(to_unsigned( 206,8)),
			13161 => std_logic_vector(to_unsigned( 219,8)),
			13162 => std_logic_vector(to_unsigned( 236,8)),
			13163 => std_logic_vector(to_unsigned( 242,8)),
			13164 => std_logic_vector(to_unsigned( 27,8)),
			13165 => std_logic_vector(to_unsigned( 4,8)),
			13166 => std_logic_vector(to_unsigned( 103,8)),
			13167 => std_logic_vector(to_unsigned( 27,8)),
			13168 => std_logic_vector(to_unsigned( 5,8)),
			13169 => std_logic_vector(to_unsigned( 239,8)),
			13170 => std_logic_vector(to_unsigned( 9,8)),
			13171 => std_logic_vector(to_unsigned( 181,8)),
			13172 => std_logic_vector(to_unsigned( 171,8)),
			13173 => std_logic_vector(to_unsigned( 171,8)),
			13174 => std_logic_vector(to_unsigned( 137,8)),
			13175 => std_logic_vector(to_unsigned( 255,8)),
			13176 => std_logic_vector(to_unsigned( 4,8)),
			13177 => std_logic_vector(to_unsigned( 78,8)),
			13178 => std_logic_vector(to_unsigned( 106,8)),
			13179 => std_logic_vector(to_unsigned( 156,8)),
			13180 => std_logic_vector(to_unsigned( 212,8)),
			13181 => std_logic_vector(to_unsigned( 116,8)),
			13182 => std_logic_vector(to_unsigned( 17,8)),
			13183 => std_logic_vector(to_unsigned( 46,8)),
			13184 => std_logic_vector(to_unsigned( 168,8)),
			13185 => std_logic_vector(to_unsigned( 98,8)),
			13186 => std_logic_vector(to_unsigned( 96,8)),
			13187 => std_logic_vector(to_unsigned( 48,8)),
			13188 => std_logic_vector(to_unsigned( 186,8)),
			13189 => std_logic_vector(to_unsigned( 249,8)),
			13190 => std_logic_vector(to_unsigned( 219,8)),
			13191 => std_logic_vector(to_unsigned( 192,8)),
			13192 => std_logic_vector(to_unsigned( 250,8)),
			13193 => std_logic_vector(to_unsigned( 29,8)),
			13194 => std_logic_vector(to_unsigned( 13,8)),
			13195 => std_logic_vector(to_unsigned( 239,8)),
			13196 => std_logic_vector(to_unsigned( 15,8)),
			13197 => std_logic_vector(to_unsigned( 75,8)),
			13198 => std_logic_vector(to_unsigned( 134,8)),
			13199 => std_logic_vector(to_unsigned( 77,8)),
			13200 => std_logic_vector(to_unsigned( 60,8)),
			13201 => std_logic_vector(to_unsigned( 203,8)),
			13202 => std_logic_vector(to_unsigned( 181,8)),
			13203 => std_logic_vector(to_unsigned( 68,8)),
			13204 => std_logic_vector(to_unsigned( 130,8)),
			13205 => std_logic_vector(to_unsigned( 2,8)),
			13206 => std_logic_vector(to_unsigned( 63,8)),
			13207 => std_logic_vector(to_unsigned( 43,8)),
			13208 => std_logic_vector(to_unsigned( 80,8)),
			13209 => std_logic_vector(to_unsigned( 144,8)),
			13210 => std_logic_vector(to_unsigned( 218,8)),
			13211 => std_logic_vector(to_unsigned( 96,8)),
			13212 => std_logic_vector(to_unsigned( 169,8)),
			13213 => std_logic_vector(to_unsigned( 183,8)),
			13214 => std_logic_vector(to_unsigned( 55,8)),
			13215 => std_logic_vector(to_unsigned( 107,8)),
			13216 => std_logic_vector(to_unsigned( 250,8)),
			13217 => std_logic_vector(to_unsigned( 60,8)),
			13218 => std_logic_vector(to_unsigned( 13,8)),
			13219 => std_logic_vector(to_unsigned( 177,8)),
			13220 => std_logic_vector(to_unsigned( 93,8)),
			13221 => std_logic_vector(to_unsigned( 221,8)),
			13222 => std_logic_vector(to_unsigned( 18,8)),
			13223 => std_logic_vector(to_unsigned( 154,8)),
			13224 => std_logic_vector(to_unsigned( 99,8)),
			13225 => std_logic_vector(to_unsigned( 243,8)),
			13226 => std_logic_vector(to_unsigned( 131,8)),
			13227 => std_logic_vector(to_unsigned( 185,8)),
			13228 => std_logic_vector(to_unsigned( 183,8)),
			13229 => std_logic_vector(to_unsigned( 224,8)),
			13230 => std_logic_vector(to_unsigned( 233,8)),
			13231 => std_logic_vector(to_unsigned( 206,8)),
			13232 => std_logic_vector(to_unsigned( 178,8)),
			13233 => std_logic_vector(to_unsigned( 195,8)),
			13234 => std_logic_vector(to_unsigned( 19,8)),
			13235 => std_logic_vector(to_unsigned( 74,8)),
			13236 => std_logic_vector(to_unsigned( 33,8)),
			13237 => std_logic_vector(to_unsigned( 40,8)),
			13238 => std_logic_vector(to_unsigned( 253,8)),
			13239 => std_logic_vector(to_unsigned( 227,8)),
			13240 => std_logic_vector(to_unsigned( 80,8)),
			13241 => std_logic_vector(to_unsigned( 51,8)),
			13242 => std_logic_vector(to_unsigned( 82,8)),
			13243 => std_logic_vector(to_unsigned( 234,8)),
			13244 => std_logic_vector(to_unsigned( 75,8)),
			13245 => std_logic_vector(to_unsigned( 120,8)),
			13246 => std_logic_vector(to_unsigned( 116,8)),
			13247 => std_logic_vector(to_unsigned( 228,8)),
			13248 => std_logic_vector(to_unsigned( 24,8)),
			13249 => std_logic_vector(to_unsigned( 13,8)),
			13250 => std_logic_vector(to_unsigned( 216,8)),
			13251 => std_logic_vector(to_unsigned( 61,8)),
			13252 => std_logic_vector(to_unsigned( 1,8)),
			13253 => std_logic_vector(to_unsigned( 59,8)),
			13254 => std_logic_vector(to_unsigned( 21,8)),
			13255 => std_logic_vector(to_unsigned( 117,8)),
			13256 => std_logic_vector(to_unsigned( 156,8)),
			13257 => std_logic_vector(to_unsigned( 254,8)),
			13258 => std_logic_vector(to_unsigned( 220,8)),
			13259 => std_logic_vector(to_unsigned( 146,8)),
			13260 => std_logic_vector(to_unsigned( 180,8)),
			13261 => std_logic_vector(to_unsigned( 145,8)),
			13262 => std_logic_vector(to_unsigned( 111,8)),
			13263 => std_logic_vector(to_unsigned( 45,8)),
			13264 => std_logic_vector(to_unsigned( 78,8)),
			13265 => std_logic_vector(to_unsigned( 19,8)),
			13266 => std_logic_vector(to_unsigned( 171,8)),
			13267 => std_logic_vector(to_unsigned( 202,8)),
			13268 => std_logic_vector(to_unsigned( 13,8)),
			13269 => std_logic_vector(to_unsigned( 72,8)),
			13270 => std_logic_vector(to_unsigned( 32,8)),
			13271 => std_logic_vector(to_unsigned( 110,8)),
			13272 => std_logic_vector(to_unsigned( 131,8)),
			13273 => std_logic_vector(to_unsigned( 153,8)),
			13274 => std_logic_vector(to_unsigned( 169,8)),
			13275 => std_logic_vector(to_unsigned( 169,8)),
			13276 => std_logic_vector(to_unsigned( 233,8)),
			13277 => std_logic_vector(to_unsigned( 176,8)),
			13278 => std_logic_vector(to_unsigned( 230,8)),
			13279 => std_logic_vector(to_unsigned( 214,8)),
			13280 => std_logic_vector(to_unsigned( 88,8)),
			13281 => std_logic_vector(to_unsigned( 103,8)),
			13282 => std_logic_vector(to_unsigned( 11,8)),
			13283 => std_logic_vector(to_unsigned( 246,8)),
			13284 => std_logic_vector(to_unsigned( 166,8)),
			13285 => std_logic_vector(to_unsigned( 96,8)),
			13286 => std_logic_vector(to_unsigned( 234,8)),
			13287 => std_logic_vector(to_unsigned( 19,8)),
			13288 => std_logic_vector(to_unsigned( 242,8)),
			13289 => std_logic_vector(to_unsigned( 35,8)),
			13290 => std_logic_vector(to_unsigned( 69,8)),
			13291 => std_logic_vector(to_unsigned( 124,8)),
			13292 => std_logic_vector(to_unsigned( 190,8)),
			13293 => std_logic_vector(to_unsigned( 158,8)),
			13294 => std_logic_vector(to_unsigned( 105,8)),
			13295 => std_logic_vector(to_unsigned( 238,8)),
			13296 => std_logic_vector(to_unsigned( 19,8)),
			13297 => std_logic_vector(to_unsigned( 45,8)),
			13298 => std_logic_vector(to_unsigned( 22,8)),
			13299 => std_logic_vector(to_unsigned( 110,8)),
			13300 => std_logic_vector(to_unsigned( 204,8)),
			13301 => std_logic_vector(to_unsigned( 75,8)),
			13302 => std_logic_vector(to_unsigned( 50,8)),
			13303 => std_logic_vector(to_unsigned( 136,8)),
			13304 => std_logic_vector(to_unsigned( 237,8)),
			13305 => std_logic_vector(to_unsigned( 17,8)),
			13306 => std_logic_vector(to_unsigned( 136,8)),
			13307 => std_logic_vector(to_unsigned( 160,8)),
			13308 => std_logic_vector(to_unsigned( 156,8)),
			13309 => std_logic_vector(to_unsigned( 8,8)),
			13310 => std_logic_vector(to_unsigned( 121,8)),
			13311 => std_logic_vector(to_unsigned( 120,8)),
			13312 => std_logic_vector(to_unsigned( 50,8)),
			13313 => std_logic_vector(to_unsigned( 247,8)),
			13314 => std_logic_vector(to_unsigned( 69,8)),
			13315 => std_logic_vector(to_unsigned( 119,8)),
			13316 => std_logic_vector(to_unsigned( 155,8)),
			13317 => std_logic_vector(to_unsigned( 194,8)),
			13318 => std_logic_vector(to_unsigned( 239,8)),
			13319 => std_logic_vector(to_unsigned( 193,8)),
			13320 => std_logic_vector(to_unsigned( 215,8)),
			13321 => std_logic_vector(to_unsigned( 45,8)),
			13322 => std_logic_vector(to_unsigned( 103,8)),
			13323 => std_logic_vector(to_unsigned( 205,8)),
			13324 => std_logic_vector(to_unsigned( 246,8)),
			13325 => std_logic_vector(to_unsigned( 242,8)),
			13326 => std_logic_vector(to_unsigned( 140,8)),
			13327 => std_logic_vector(to_unsigned( 214,8)),
			13328 => std_logic_vector(to_unsigned( 38,8)),
			13329 => std_logic_vector(to_unsigned( 55,8)),
			13330 => std_logic_vector(to_unsigned( 147,8)),
			13331 => std_logic_vector(to_unsigned( 59,8)),
			13332 => std_logic_vector(to_unsigned( 124,8)),
			13333 => std_logic_vector(to_unsigned( 114,8)),
			13334 => std_logic_vector(to_unsigned( 241,8)),
			13335 => std_logic_vector(to_unsigned( 163,8)),
			13336 => std_logic_vector(to_unsigned( 20,8)),
			13337 => std_logic_vector(to_unsigned( 49,8)),
			13338 => std_logic_vector(to_unsigned( 122,8)),
			13339 => std_logic_vector(to_unsigned( 193,8)),
			13340 => std_logic_vector(to_unsigned( 180,8)),
			13341 => std_logic_vector(to_unsigned( 105,8)),
			13342 => std_logic_vector(to_unsigned( 137,8)),
			13343 => std_logic_vector(to_unsigned( 177,8)),
			13344 => std_logic_vector(to_unsigned( 181,8)),
			13345 => std_logic_vector(to_unsigned( 122,8)),
			13346 => std_logic_vector(to_unsigned( 130,8)),
			13347 => std_logic_vector(to_unsigned( 76,8)),
			13348 => std_logic_vector(to_unsigned( 232,8)),
			13349 => std_logic_vector(to_unsigned( 226,8)),
			13350 => std_logic_vector(to_unsigned( 29,8)),
			13351 => std_logic_vector(to_unsigned( 38,8)),
			13352 => std_logic_vector(to_unsigned( 32,8)),
			13353 => std_logic_vector(to_unsigned( 133,8)),
			13354 => std_logic_vector(to_unsigned( 57,8)),
			13355 => std_logic_vector(to_unsigned( 126,8)),
			13356 => std_logic_vector(to_unsigned( 168,8)),
			13357 => std_logic_vector(to_unsigned( 121,8)),
			13358 => std_logic_vector(to_unsigned( 27,8)),
			13359 => std_logic_vector(to_unsigned( 10,8)),
			13360 => std_logic_vector(to_unsigned( 52,8)),
			13361 => std_logic_vector(to_unsigned( 210,8)),
			13362 => std_logic_vector(to_unsigned( 236,8)),
			13363 => std_logic_vector(to_unsigned( 14,8)),
			13364 => std_logic_vector(to_unsigned( 175,8)),
			13365 => std_logic_vector(to_unsigned( 50,8)),
			13366 => std_logic_vector(to_unsigned( 204,8)),
			13367 => std_logic_vector(to_unsigned( 70,8)),
			13368 => std_logic_vector(to_unsigned( 240,8)),
			13369 => std_logic_vector(to_unsigned( 68,8)),
			13370 => std_logic_vector(to_unsigned( 103,8)),
			13371 => std_logic_vector(to_unsigned( 239,8)),
			13372 => std_logic_vector(to_unsigned( 4,8)),
			13373 => std_logic_vector(to_unsigned( 47,8)),
			13374 => std_logic_vector(to_unsigned( 8,8)),
			13375 => std_logic_vector(to_unsigned( 112,8)),
			13376 => std_logic_vector(to_unsigned( 43,8)),
			13377 => std_logic_vector(to_unsigned( 174,8)),
			13378 => std_logic_vector(to_unsigned( 96,8)),
			13379 => std_logic_vector(to_unsigned( 156,8)),
			13380 => std_logic_vector(to_unsigned( 74,8)),
			13381 => std_logic_vector(to_unsigned( 235,8)),
			13382 => std_logic_vector(to_unsigned( 13,8)),
			13383 => std_logic_vector(to_unsigned( 1,8)),
			13384 => std_logic_vector(to_unsigned( 71,8)),
			13385 => std_logic_vector(to_unsigned( 37,8)),
			13386 => std_logic_vector(to_unsigned( 220,8)),
			13387 => std_logic_vector(to_unsigned( 153,8)),
			13388 => std_logic_vector(to_unsigned( 109,8)),
			13389 => std_logic_vector(to_unsigned( 213,8)),
			13390 => std_logic_vector(to_unsigned( 117,8)),
			13391 => std_logic_vector(to_unsigned( 80,8)),
			13392 => std_logic_vector(to_unsigned( 39,8)),
			13393 => std_logic_vector(to_unsigned( 51,8)),
			13394 => std_logic_vector(to_unsigned( 249,8)),
			13395 => std_logic_vector(to_unsigned( 7,8)),
			13396 => std_logic_vector(to_unsigned( 253,8)),
			13397 => std_logic_vector(to_unsigned( 175,8)),
			13398 => std_logic_vector(to_unsigned( 45,8)),
			13399 => std_logic_vector(to_unsigned( 195,8)),
			13400 => std_logic_vector(to_unsigned( 141,8)),
			13401 => std_logic_vector(to_unsigned( 98,8)),
			13402 => std_logic_vector(to_unsigned( 188,8)),
			13403 => std_logic_vector(to_unsigned( 34,8)),
			13404 => std_logic_vector(to_unsigned( 168,8)),
			13405 => std_logic_vector(to_unsigned( 169,8)),
			13406 => std_logic_vector(to_unsigned( 133,8)),
			13407 => std_logic_vector(to_unsigned( 243,8)),
			13408 => std_logic_vector(to_unsigned( 238,8)),
			13409 => std_logic_vector(to_unsigned( 33,8)),
			13410 => std_logic_vector(to_unsigned( 21,8)),
			13411 => std_logic_vector(to_unsigned( 213,8)),
			13412 => std_logic_vector(to_unsigned( 225,8)),
			13413 => std_logic_vector(to_unsigned( 119,8)),
			13414 => std_logic_vector(to_unsigned( 141,8)),
			13415 => std_logic_vector(to_unsigned( 120,8)),
			13416 => std_logic_vector(to_unsigned( 101,8)),
			13417 => std_logic_vector(to_unsigned( 73,8)),
			13418 => std_logic_vector(to_unsigned( 146,8)),
			13419 => std_logic_vector(to_unsigned( 141,8)),
			13420 => std_logic_vector(to_unsigned( 126,8)),
			13421 => std_logic_vector(to_unsigned( 129,8)),
			13422 => std_logic_vector(to_unsigned( 213,8)),
			13423 => std_logic_vector(to_unsigned( 80,8)),
			13424 => std_logic_vector(to_unsigned( 152,8)),
			13425 => std_logic_vector(to_unsigned( 63,8)),
			13426 => std_logic_vector(to_unsigned( 94,8)),
			13427 => std_logic_vector(to_unsigned( 116,8)),
			13428 => std_logic_vector(to_unsigned( 15,8)),
			13429 => std_logic_vector(to_unsigned( 26,8)),
			13430 => std_logic_vector(to_unsigned( 7,8)),
			13431 => std_logic_vector(to_unsigned( 204,8)),
			13432 => std_logic_vector(to_unsigned( 255,8)),
			13433 => std_logic_vector(to_unsigned( 63,8)),
			13434 => std_logic_vector(to_unsigned( 125,8)),
			13435 => std_logic_vector(to_unsigned( 204,8)),
			13436 => std_logic_vector(to_unsigned( 81,8)),
			13437 => std_logic_vector(to_unsigned( 204,8)),
			13438 => std_logic_vector(to_unsigned( 69,8)),
			13439 => std_logic_vector(to_unsigned( 134,8)),
			13440 => std_logic_vector(to_unsigned( 147,8)),
			13441 => std_logic_vector(to_unsigned( 217,8)),
			13442 => std_logic_vector(to_unsigned( 86,8)),
			13443 => std_logic_vector(to_unsigned( 124,8)),
			13444 => std_logic_vector(to_unsigned( 120,8)),
			13445 => std_logic_vector(to_unsigned( 7,8)),
			13446 => std_logic_vector(to_unsigned( 26,8)),
			13447 => std_logic_vector(to_unsigned( 87,8)),
			13448 => std_logic_vector(to_unsigned( 130,8)),
			13449 => std_logic_vector(to_unsigned( 248,8)),
			13450 => std_logic_vector(to_unsigned( 207,8)),
			13451 => std_logic_vector(to_unsigned( 146,8)),
			13452 => std_logic_vector(to_unsigned( 132,8)),
			13453 => std_logic_vector(to_unsigned( 22,8)),
			13454 => std_logic_vector(to_unsigned( 2,8)),
			13455 => std_logic_vector(to_unsigned( 49,8)),
			13456 => std_logic_vector(to_unsigned( 109,8)),
			13457 => std_logic_vector(to_unsigned( 44,8)),
			13458 => std_logic_vector(to_unsigned( 228,8)),
			13459 => std_logic_vector(to_unsigned( 181,8)),
			13460 => std_logic_vector(to_unsigned( 164,8)),
			13461 => std_logic_vector(to_unsigned( 18,8)),
			13462 => std_logic_vector(to_unsigned( 22,8)),
			13463 => std_logic_vector(to_unsigned( 188,8)),
			13464 => std_logic_vector(to_unsigned( 123,8)),
			13465 => std_logic_vector(to_unsigned( 80,8)),
			13466 => std_logic_vector(to_unsigned( 163,8)),
			13467 => std_logic_vector(to_unsigned( 9,8)),
			13468 => std_logic_vector(to_unsigned( 85,8)),
			13469 => std_logic_vector(to_unsigned( 239,8)),
			13470 => std_logic_vector(to_unsigned( 142,8)),
			13471 => std_logic_vector(to_unsigned( 176,8)),
			13472 => std_logic_vector(to_unsigned( 202,8)),
			13473 => std_logic_vector(to_unsigned( 25,8)),
			13474 => std_logic_vector(to_unsigned( 93,8)),
			13475 => std_logic_vector(to_unsigned( 71,8)),
			13476 => std_logic_vector(to_unsigned( 25,8)),
			13477 => std_logic_vector(to_unsigned( 211,8)),
			13478 => std_logic_vector(to_unsigned( 67,8)),
			13479 => std_logic_vector(to_unsigned( 85,8)),
			13480 => std_logic_vector(to_unsigned( 228,8)),
			13481 => std_logic_vector(to_unsigned( 252,8)),
			13482 => std_logic_vector(to_unsigned( 81,8)),
			13483 => std_logic_vector(to_unsigned( 248,8)),
			13484 => std_logic_vector(to_unsigned( 156,8)),
			13485 => std_logic_vector(to_unsigned( 171,8)),
			13486 => std_logic_vector(to_unsigned( 40,8)),
			13487 => std_logic_vector(to_unsigned( 164,8)),
			13488 => std_logic_vector(to_unsigned( 203,8)),
			13489 => std_logic_vector(to_unsigned( 208,8)),
			13490 => std_logic_vector(to_unsigned( 212,8)),
			13491 => std_logic_vector(to_unsigned( 249,8)),
			13492 => std_logic_vector(to_unsigned( 111,8)),
			13493 => std_logic_vector(to_unsigned( 46,8)),
			13494 => std_logic_vector(to_unsigned( 167,8)),
			13495 => std_logic_vector(to_unsigned( 139,8)),
			13496 => std_logic_vector(to_unsigned( 39,8)),
			13497 => std_logic_vector(to_unsigned( 146,8)),
			13498 => std_logic_vector(to_unsigned( 149,8)),
			13499 => std_logic_vector(to_unsigned( 167,8)),
			13500 => std_logic_vector(to_unsigned( 228,8)),
			13501 => std_logic_vector(to_unsigned( 173,8)),
			13502 => std_logic_vector(to_unsigned( 5,8)),
			13503 => std_logic_vector(to_unsigned( 151,8)),
			13504 => std_logic_vector(to_unsigned( 150,8)),
			13505 => std_logic_vector(to_unsigned( 158,8)),
			13506 => std_logic_vector(to_unsigned( 253,8)),
			13507 => std_logic_vector(to_unsigned( 56,8)),
			13508 => std_logic_vector(to_unsigned( 230,8)),
			13509 => std_logic_vector(to_unsigned( 138,8)),
			13510 => std_logic_vector(to_unsigned( 70,8)),
			13511 => std_logic_vector(to_unsigned( 230,8)),
			13512 => std_logic_vector(to_unsigned( 23,8)),
			13513 => std_logic_vector(to_unsigned( 17,8)),
			13514 => std_logic_vector(to_unsigned( 167,8)),
			13515 => std_logic_vector(to_unsigned( 112,8)),
			13516 => std_logic_vector(to_unsigned( 152,8)),
			13517 => std_logic_vector(to_unsigned( 90,8)),
			13518 => std_logic_vector(to_unsigned( 68,8)),
			13519 => std_logic_vector(to_unsigned( 20,8)),
			13520 => std_logic_vector(to_unsigned( 15,8)),
			13521 => std_logic_vector(to_unsigned( 10,8)),
			13522 => std_logic_vector(to_unsigned( 125,8)),
			13523 => std_logic_vector(to_unsigned( 247,8)),
			13524 => std_logic_vector(to_unsigned( 200,8)),
			13525 => std_logic_vector(to_unsigned( 108,8)),
			13526 => std_logic_vector(to_unsigned( 157,8)),
			13527 => std_logic_vector(to_unsigned( 30,8)),
			13528 => std_logic_vector(to_unsigned( 21,8)),
			13529 => std_logic_vector(to_unsigned( 249,8)),
			13530 => std_logic_vector(to_unsigned( 202,8)),
			13531 => std_logic_vector(to_unsigned( 6,8)),
			13532 => std_logic_vector(to_unsigned( 147,8)),
			13533 => std_logic_vector(to_unsigned( 34,8)),
			13534 => std_logic_vector(to_unsigned( 29,8)),
			13535 => std_logic_vector(to_unsigned( 194,8)),
			13536 => std_logic_vector(to_unsigned( 77,8)),
			13537 => std_logic_vector(to_unsigned( 224,8)),
			13538 => std_logic_vector(to_unsigned( 116,8)),
			13539 => std_logic_vector(to_unsigned( 84,8)),
			13540 => std_logic_vector(to_unsigned( 177,8)),
			13541 => std_logic_vector(to_unsigned( 111,8)),
			13542 => std_logic_vector(to_unsigned( 59,8)),
			13543 => std_logic_vector(to_unsigned( 119,8)),
			13544 => std_logic_vector(to_unsigned( 145,8)),
			13545 => std_logic_vector(to_unsigned( 94,8)),
			13546 => std_logic_vector(to_unsigned( 57,8)),
			13547 => std_logic_vector(to_unsigned( 113,8)),
			13548 => std_logic_vector(to_unsigned( 8,8)),
			13549 => std_logic_vector(to_unsigned( 144,8)),
			13550 => std_logic_vector(to_unsigned( 11,8)),
			13551 => std_logic_vector(to_unsigned( 106,8)),
			13552 => std_logic_vector(to_unsigned( 10,8)),
			13553 => std_logic_vector(to_unsigned( 76,8)),
			13554 => std_logic_vector(to_unsigned( 146,8)),
			13555 => std_logic_vector(to_unsigned( 191,8)),
			13556 => std_logic_vector(to_unsigned( 128,8)),
			13557 => std_logic_vector(to_unsigned( 153,8)),
			13558 => std_logic_vector(to_unsigned( 238,8)),
			13559 => std_logic_vector(to_unsigned( 163,8)),
			13560 => std_logic_vector(to_unsigned( 178,8)),
			13561 => std_logic_vector(to_unsigned( 212,8)),
			13562 => std_logic_vector(to_unsigned( 133,8)),
			13563 => std_logic_vector(to_unsigned( 228,8)),
			13564 => std_logic_vector(to_unsigned( 185,8)),
			13565 => std_logic_vector(to_unsigned( 30,8)),
			13566 => std_logic_vector(to_unsigned( 88,8)),
			13567 => std_logic_vector(to_unsigned( 198,8)),
			13568 => std_logic_vector(to_unsigned( 214,8)),
			13569 => std_logic_vector(to_unsigned( 193,8)),
			13570 => std_logic_vector(to_unsigned( 0,8)),
			13571 => std_logic_vector(to_unsigned( 169,8)),
			13572 => std_logic_vector(to_unsigned( 136,8)),
			13573 => std_logic_vector(to_unsigned( 221,8)),
			13574 => std_logic_vector(to_unsigned( 75,8)),
			13575 => std_logic_vector(to_unsigned( 72,8)),
			13576 => std_logic_vector(to_unsigned( 52,8)),
			13577 => std_logic_vector(to_unsigned( 163,8)),
			13578 => std_logic_vector(to_unsigned( 198,8)),
			13579 => std_logic_vector(to_unsigned( 76,8)),
			13580 => std_logic_vector(to_unsigned( 32,8)),
			13581 => std_logic_vector(to_unsigned( 142,8)),
			13582 => std_logic_vector(to_unsigned( 166,8)),
			13583 => std_logic_vector(to_unsigned( 61,8)),
			13584 => std_logic_vector(to_unsigned( 12,8)),
			13585 => std_logic_vector(to_unsigned( 190,8)),
			13586 => std_logic_vector(to_unsigned( 98,8)),
			13587 => std_logic_vector(to_unsigned( 61,8)),
			13588 => std_logic_vector(to_unsigned( 117,8)),
			13589 => std_logic_vector(to_unsigned( 145,8)),
			13590 => std_logic_vector(to_unsigned( 181,8)),
			13591 => std_logic_vector(to_unsigned( 193,8)),
			13592 => std_logic_vector(to_unsigned( 197,8)),
			13593 => std_logic_vector(to_unsigned( 247,8)),
			13594 => std_logic_vector(to_unsigned( 171,8)),
			13595 => std_logic_vector(to_unsigned( 27,8)),
			13596 => std_logic_vector(to_unsigned( 180,8)),
			13597 => std_logic_vector(to_unsigned( 111,8)),
			13598 => std_logic_vector(to_unsigned( 193,8)),
			13599 => std_logic_vector(to_unsigned( 139,8)),
			13600 => std_logic_vector(to_unsigned( 147,8)),
			13601 => std_logic_vector(to_unsigned( 187,8)),
			13602 => std_logic_vector(to_unsigned( 17,8)),
			13603 => std_logic_vector(to_unsigned( 230,8)),
			13604 => std_logic_vector(to_unsigned( 44,8)),
			13605 => std_logic_vector(to_unsigned( 106,8)),
			13606 => std_logic_vector(to_unsigned( 6,8)),
			13607 => std_logic_vector(to_unsigned( 91,8)),
			13608 => std_logic_vector(to_unsigned( 62,8)),
			13609 => std_logic_vector(to_unsigned( 230,8)),
			13610 => std_logic_vector(to_unsigned( 15,8)),
			13611 => std_logic_vector(to_unsigned( 118,8)),
			13612 => std_logic_vector(to_unsigned( 172,8)),
			13613 => std_logic_vector(to_unsigned( 119,8)),
			13614 => std_logic_vector(to_unsigned( 119,8)),
			13615 => std_logic_vector(to_unsigned( 154,8)),
			13616 => std_logic_vector(to_unsigned( 164,8)),
			13617 => std_logic_vector(to_unsigned( 13,8)),
			13618 => std_logic_vector(to_unsigned( 168,8)),
			13619 => std_logic_vector(to_unsigned( 159,8)),
			13620 => std_logic_vector(to_unsigned( 55,8)),
			13621 => std_logic_vector(to_unsigned( 139,8)),
			13622 => std_logic_vector(to_unsigned( 47,8)),
			13623 => std_logic_vector(to_unsigned( 176,8)),
			13624 => std_logic_vector(to_unsigned( 194,8)),
			13625 => std_logic_vector(to_unsigned( 51,8)),
			13626 => std_logic_vector(to_unsigned( 126,8)),
			13627 => std_logic_vector(to_unsigned( 78,8)),
			13628 => std_logic_vector(to_unsigned( 92,8)),
			13629 => std_logic_vector(to_unsigned( 40,8)),
			13630 => std_logic_vector(to_unsigned( 148,8)),
			13631 => std_logic_vector(to_unsigned( 27,8)),
			13632 => std_logic_vector(to_unsigned( 136,8)),
			13633 => std_logic_vector(to_unsigned( 219,8)),
			13634 => std_logic_vector(to_unsigned( 223,8)),
			13635 => std_logic_vector(to_unsigned( 169,8)),
			13636 => std_logic_vector(to_unsigned( 21,8)),
			13637 => std_logic_vector(to_unsigned( 205,8)),
			13638 => std_logic_vector(to_unsigned( 48,8)),
			13639 => std_logic_vector(to_unsigned( 206,8)),
			13640 => std_logic_vector(to_unsigned( 15,8)),
			13641 => std_logic_vector(to_unsigned( 195,8)),
			13642 => std_logic_vector(to_unsigned( 247,8)),
			13643 => std_logic_vector(to_unsigned( 178,8)),
			13644 => std_logic_vector(to_unsigned( 235,8)),
			13645 => std_logic_vector(to_unsigned( 179,8)),
			13646 => std_logic_vector(to_unsigned( 151,8)),
			13647 => std_logic_vector(to_unsigned( 95,8)),
			13648 => std_logic_vector(to_unsigned( 166,8)),
			13649 => std_logic_vector(to_unsigned( 45,8)),
			13650 => std_logic_vector(to_unsigned( 233,8)),
			13651 => std_logic_vector(to_unsigned( 193,8)),
			13652 => std_logic_vector(to_unsigned( 184,8)),
			13653 => std_logic_vector(to_unsigned( 234,8)),
			13654 => std_logic_vector(to_unsigned( 61,8)),
			13655 => std_logic_vector(to_unsigned( 2,8)),
			13656 => std_logic_vector(to_unsigned( 3,8)),
			13657 => std_logic_vector(to_unsigned( 51,8)),
			13658 => std_logic_vector(to_unsigned( 178,8)),
			13659 => std_logic_vector(to_unsigned( 165,8)),
			13660 => std_logic_vector(to_unsigned( 45,8)),
			13661 => std_logic_vector(to_unsigned( 40,8)),
			13662 => std_logic_vector(to_unsigned( 154,8)),
			13663 => std_logic_vector(to_unsigned( 11,8)),
			13664 => std_logic_vector(to_unsigned( 49,8)),
			13665 => std_logic_vector(to_unsigned( 205,8)),
			13666 => std_logic_vector(to_unsigned( 17,8)),
			13667 => std_logic_vector(to_unsigned( 152,8)),
			13668 => std_logic_vector(to_unsigned( 66,8)),
			13669 => std_logic_vector(to_unsigned( 194,8)),
			13670 => std_logic_vector(to_unsigned( 209,8)),
			13671 => std_logic_vector(to_unsigned( 49,8)),
			13672 => std_logic_vector(to_unsigned( 228,8)),
			13673 => std_logic_vector(to_unsigned( 133,8)),
			13674 => std_logic_vector(to_unsigned( 177,8)),
			13675 => std_logic_vector(to_unsigned( 223,8)),
			13676 => std_logic_vector(to_unsigned( 236,8)),
			13677 => std_logic_vector(to_unsigned( 198,8)),
			13678 => std_logic_vector(to_unsigned( 105,8)),
			13679 => std_logic_vector(to_unsigned( 112,8)),
			13680 => std_logic_vector(to_unsigned( 116,8)),
			13681 => std_logic_vector(to_unsigned( 117,8)),
			13682 => std_logic_vector(to_unsigned( 206,8)),
			13683 => std_logic_vector(to_unsigned( 58,8)),
			13684 => std_logic_vector(to_unsigned( 37,8)),
			13685 => std_logic_vector(to_unsigned( 116,8)),
			13686 => std_logic_vector(to_unsigned( 3,8)),
			13687 => std_logic_vector(to_unsigned( 57,8)),
			13688 => std_logic_vector(to_unsigned( 43,8)),
			13689 => std_logic_vector(to_unsigned( 185,8)),
			13690 => std_logic_vector(to_unsigned( 172,8)),
			13691 => std_logic_vector(to_unsigned( 227,8)),
			13692 => std_logic_vector(to_unsigned( 210,8)),
			13693 => std_logic_vector(to_unsigned( 78,8)),
			13694 => std_logic_vector(to_unsigned( 151,8)),
			13695 => std_logic_vector(to_unsigned( 215,8)),
			13696 => std_logic_vector(to_unsigned( 199,8)),
			13697 => std_logic_vector(to_unsigned( 234,8)),
			13698 => std_logic_vector(to_unsigned( 119,8)),
			13699 => std_logic_vector(to_unsigned( 176,8)),
			13700 => std_logic_vector(to_unsigned( 71,8)),
			13701 => std_logic_vector(to_unsigned( 241,8)),
			13702 => std_logic_vector(to_unsigned( 31,8)),
			13703 => std_logic_vector(to_unsigned( 62,8)),
			13704 => std_logic_vector(to_unsigned( 210,8)),
			13705 => std_logic_vector(to_unsigned( 215,8)),
			13706 => std_logic_vector(to_unsigned( 21,8)),
			13707 => std_logic_vector(to_unsigned( 137,8)),
			13708 => std_logic_vector(to_unsigned( 58,8)),
			13709 => std_logic_vector(to_unsigned( 243,8)),
			13710 => std_logic_vector(to_unsigned( 13,8)),
			13711 => std_logic_vector(to_unsigned( 30,8)),
			13712 => std_logic_vector(to_unsigned( 163,8)),
			13713 => std_logic_vector(to_unsigned( 126,8)),
			13714 => std_logic_vector(to_unsigned( 235,8)),
			13715 => std_logic_vector(to_unsigned( 127,8)),
			13716 => std_logic_vector(to_unsigned( 111,8)),
			13717 => std_logic_vector(to_unsigned( 187,8)),
			13718 => std_logic_vector(to_unsigned( 146,8)),
			13719 => std_logic_vector(to_unsigned( 58,8)),
			13720 => std_logic_vector(to_unsigned( 67,8)),
			13721 => std_logic_vector(to_unsigned( 7,8)),
			13722 => std_logic_vector(to_unsigned( 3,8)),
			13723 => std_logic_vector(to_unsigned( 28,8)),
			13724 => std_logic_vector(to_unsigned( 232,8)),
			13725 => std_logic_vector(to_unsigned( 3,8)),
			13726 => std_logic_vector(to_unsigned( 31,8)),
			13727 => std_logic_vector(to_unsigned( 4,8)),
			13728 => std_logic_vector(to_unsigned( 161,8)),
			13729 => std_logic_vector(to_unsigned( 254,8)),
			13730 => std_logic_vector(to_unsigned( 42,8)),
			13731 => std_logic_vector(to_unsigned( 125,8)),
			13732 => std_logic_vector(to_unsigned( 157,8)),
			13733 => std_logic_vector(to_unsigned( 161,8)),
			13734 => std_logic_vector(to_unsigned( 5,8)),
			13735 => std_logic_vector(to_unsigned( 38,8)),
			13736 => std_logic_vector(to_unsigned( 161,8)),
			13737 => std_logic_vector(to_unsigned( 97,8)),
			13738 => std_logic_vector(to_unsigned( 228,8)),
			13739 => std_logic_vector(to_unsigned( 250,8)),
			13740 => std_logic_vector(to_unsigned( 136,8)),
			13741 => std_logic_vector(to_unsigned( 4,8)),
			13742 => std_logic_vector(to_unsigned( 42,8)),
			13743 => std_logic_vector(to_unsigned( 173,8)),
			13744 => std_logic_vector(to_unsigned( 91,8)),
			13745 => std_logic_vector(to_unsigned( 122,8)),
			13746 => std_logic_vector(to_unsigned( 79,8)),
			13747 => std_logic_vector(to_unsigned( 34,8)),
			13748 => std_logic_vector(to_unsigned( 204,8)),
			13749 => std_logic_vector(to_unsigned( 196,8)),
			13750 => std_logic_vector(to_unsigned( 133,8)),
			13751 => std_logic_vector(to_unsigned( 238,8)),
			13752 => std_logic_vector(to_unsigned( 17,8)),
			13753 => std_logic_vector(to_unsigned( 122,8)),
			13754 => std_logic_vector(to_unsigned( 73,8)),
			13755 => std_logic_vector(to_unsigned( 225,8)),
			13756 => std_logic_vector(to_unsigned( 186,8)),
			13757 => std_logic_vector(to_unsigned( 103,8)),
			13758 => std_logic_vector(to_unsigned( 185,8)),
			13759 => std_logic_vector(to_unsigned( 146,8)),
			13760 => std_logic_vector(to_unsigned( 193,8)),
			13761 => std_logic_vector(to_unsigned( 238,8)),
			13762 => std_logic_vector(to_unsigned( 75,8)),
			13763 => std_logic_vector(to_unsigned( 11,8)),
			13764 => std_logic_vector(to_unsigned( 120,8)),
			13765 => std_logic_vector(to_unsigned( 207,8)),
			13766 => std_logic_vector(to_unsigned( 5,8)),
			13767 => std_logic_vector(to_unsigned( 14,8)),
			13768 => std_logic_vector(to_unsigned( 99,8)),
			13769 => std_logic_vector(to_unsigned( 75,8)),
			13770 => std_logic_vector(to_unsigned( 209,8)),
			13771 => std_logic_vector(to_unsigned( 227,8)),
			13772 => std_logic_vector(to_unsigned( 134,8)),
			13773 => std_logic_vector(to_unsigned( 28,8)),
			13774 => std_logic_vector(to_unsigned( 121,8)),
			13775 => std_logic_vector(to_unsigned( 226,8)),
			13776 => std_logic_vector(to_unsigned( 159,8)),
			13777 => std_logic_vector(to_unsigned( 231,8)),
			13778 => std_logic_vector(to_unsigned( 21,8)),
			13779 => std_logic_vector(to_unsigned( 185,8)),
			13780 => std_logic_vector(to_unsigned( 93,8)),
			13781 => std_logic_vector(to_unsigned( 133,8)),
			13782 => std_logic_vector(to_unsigned( 67,8)),
			13783 => std_logic_vector(to_unsigned( 53,8)),
			13784 => std_logic_vector(to_unsigned( 200,8)),
			13785 => std_logic_vector(to_unsigned( 206,8)),
			13786 => std_logic_vector(to_unsigned( 219,8)),
			13787 => std_logic_vector(to_unsigned( 179,8)),
			13788 => std_logic_vector(to_unsigned( 25,8)),
			13789 => std_logic_vector(to_unsigned( 202,8)),
			13790 => std_logic_vector(to_unsigned( 155,8)),
			13791 => std_logic_vector(to_unsigned( 138,8)),
			13792 => std_logic_vector(to_unsigned( 8,8)),
			13793 => std_logic_vector(to_unsigned( 160,8)),
			13794 => std_logic_vector(to_unsigned( 22,8)),
			13795 => std_logic_vector(to_unsigned( 176,8)),
			13796 => std_logic_vector(to_unsigned( 205,8)),
			13797 => std_logic_vector(to_unsigned( 39,8)),
			13798 => std_logic_vector(to_unsigned( 194,8)),
			13799 => std_logic_vector(to_unsigned( 71,8)),
			13800 => std_logic_vector(to_unsigned( 9,8)),
			13801 => std_logic_vector(to_unsigned( 31,8)),
			13802 => std_logic_vector(to_unsigned( 213,8)),
			13803 => std_logic_vector(to_unsigned( 186,8)),
			13804 => std_logic_vector(to_unsigned( 8,8)),
			13805 => std_logic_vector(to_unsigned( 176,8)),
			13806 => std_logic_vector(to_unsigned( 86,8)),
			13807 => std_logic_vector(to_unsigned( 228,8)),
			13808 => std_logic_vector(to_unsigned( 168,8)),
			13809 => std_logic_vector(to_unsigned( 219,8)),
			13810 => std_logic_vector(to_unsigned( 180,8)),
			13811 => std_logic_vector(to_unsigned( 50,8)),
			13812 => std_logic_vector(to_unsigned( 94,8)),
			13813 => std_logic_vector(to_unsigned( 83,8)),
			13814 => std_logic_vector(to_unsigned( 111,8)),
			13815 => std_logic_vector(to_unsigned( 71,8)),
			13816 => std_logic_vector(to_unsigned( 190,8)),
			13817 => std_logic_vector(to_unsigned( 15,8)),
			13818 => std_logic_vector(to_unsigned( 235,8)),
			13819 => std_logic_vector(to_unsigned( 182,8)),
			13820 => std_logic_vector(to_unsigned( 131,8)),
			13821 => std_logic_vector(to_unsigned( 98,8)),
			13822 => std_logic_vector(to_unsigned( 155,8)),
			13823 => std_logic_vector(to_unsigned( 97,8)),
			13824 => std_logic_vector(to_unsigned( 83,8)),
			13825 => std_logic_vector(to_unsigned( 193,8)),
			13826 => std_logic_vector(to_unsigned( 3,8)),
			13827 => std_logic_vector(to_unsigned( 165,8)),
			13828 => std_logic_vector(to_unsigned( 171,8)),
			13829 => std_logic_vector(to_unsigned( 195,8)),
			13830 => std_logic_vector(to_unsigned( 239,8)),
			13831 => std_logic_vector(to_unsigned( 177,8)),
			13832 => std_logic_vector(to_unsigned( 95,8)),
			13833 => std_logic_vector(to_unsigned( 67,8)),
			13834 => std_logic_vector(to_unsigned( 65,8)),
			13835 => std_logic_vector(to_unsigned( 243,8)),
			13836 => std_logic_vector(to_unsigned( 188,8)),
			13837 => std_logic_vector(to_unsigned( 107,8)),
			13838 => std_logic_vector(to_unsigned( 150,8)),
			13839 => std_logic_vector(to_unsigned( 16,8)),
			13840 => std_logic_vector(to_unsigned( 10,8)),
			13841 => std_logic_vector(to_unsigned( 201,8)),
			13842 => std_logic_vector(to_unsigned( 46,8)),
			13843 => std_logic_vector(to_unsigned( 45,8)),
			13844 => std_logic_vector(to_unsigned( 128,8)),
			13845 => std_logic_vector(to_unsigned( 139,8)),
			13846 => std_logic_vector(to_unsigned( 193,8)),
			13847 => std_logic_vector(to_unsigned( 95,8)),
			13848 => std_logic_vector(to_unsigned( 206,8)),
			13849 => std_logic_vector(to_unsigned( 72,8)),
			13850 => std_logic_vector(to_unsigned( 107,8)),
			13851 => std_logic_vector(to_unsigned( 154,8)),
			13852 => std_logic_vector(to_unsigned( 18,8)),
			13853 => std_logic_vector(to_unsigned( 74,8)),
			13854 => std_logic_vector(to_unsigned( 139,8)),
			13855 => std_logic_vector(to_unsigned( 71,8)),
			13856 => std_logic_vector(to_unsigned( 26,8)),
			13857 => std_logic_vector(to_unsigned( 51,8)),
			13858 => std_logic_vector(to_unsigned( 185,8)),
			13859 => std_logic_vector(to_unsigned( 17,8)),
			13860 => std_logic_vector(to_unsigned( 222,8)),
			13861 => std_logic_vector(to_unsigned( 214,8)),
			13862 => std_logic_vector(to_unsigned( 166,8)),
			13863 => std_logic_vector(to_unsigned( 208,8)),
			13864 => std_logic_vector(to_unsigned( 59,8)),
			13865 => std_logic_vector(to_unsigned( 125,8)),
			13866 => std_logic_vector(to_unsigned( 31,8)),
			13867 => std_logic_vector(to_unsigned( 180,8)),
			13868 => std_logic_vector(to_unsigned( 223,8)),
			13869 => std_logic_vector(to_unsigned( 52,8)),
			13870 => std_logic_vector(to_unsigned( 2,8)),
			13871 => std_logic_vector(to_unsigned( 102,8)),
			13872 => std_logic_vector(to_unsigned( 244,8)),
			13873 => std_logic_vector(to_unsigned( 164,8)),
			13874 => std_logic_vector(to_unsigned( 196,8)),
			13875 => std_logic_vector(to_unsigned( 21,8)),
			13876 => std_logic_vector(to_unsigned( 133,8)),
			13877 => std_logic_vector(to_unsigned( 227,8)),
			13878 => std_logic_vector(to_unsigned( 111,8)),
			13879 => std_logic_vector(to_unsigned( 72,8)),
			13880 => std_logic_vector(to_unsigned( 200,8)),
			13881 => std_logic_vector(to_unsigned( 4,8)),
			13882 => std_logic_vector(to_unsigned( 219,8)),
			13883 => std_logic_vector(to_unsigned( 188,8)),
			13884 => std_logic_vector(to_unsigned( 189,8)),
			13885 => std_logic_vector(to_unsigned( 25,8)),
			13886 => std_logic_vector(to_unsigned( 229,8)),
			13887 => std_logic_vector(to_unsigned( 253,8)),
			13888 => std_logic_vector(to_unsigned( 27,8)),
			13889 => std_logic_vector(to_unsigned( 229,8)),
			13890 => std_logic_vector(to_unsigned( 217,8)),
			13891 => std_logic_vector(to_unsigned( 202,8)),
			13892 => std_logic_vector(to_unsigned( 248,8)),
			13893 => std_logic_vector(to_unsigned( 13,8)),
			13894 => std_logic_vector(to_unsigned( 110,8)),
			13895 => std_logic_vector(to_unsigned( 238,8)),
			13896 => std_logic_vector(to_unsigned( 19,8)),
			13897 => std_logic_vector(to_unsigned( 192,8)),
			13898 => std_logic_vector(to_unsigned( 16,8)),
			13899 => std_logic_vector(to_unsigned( 160,8)),
			13900 => std_logic_vector(to_unsigned( 214,8)),
			13901 => std_logic_vector(to_unsigned( 221,8)),
			13902 => std_logic_vector(to_unsigned( 191,8)),
			13903 => std_logic_vector(to_unsigned( 164,8)),
			13904 => std_logic_vector(to_unsigned( 198,8)),
			13905 => std_logic_vector(to_unsigned( 83,8)),
			13906 => std_logic_vector(to_unsigned( 191,8)),
			13907 => std_logic_vector(to_unsigned( 180,8)),
			13908 => std_logic_vector(to_unsigned( 180,8)),
			13909 => std_logic_vector(to_unsigned( 113,8)),
			13910 => std_logic_vector(to_unsigned( 162,8)),
			13911 => std_logic_vector(to_unsigned( 103,8)),
			13912 => std_logic_vector(to_unsigned( 230,8)),
			13913 => std_logic_vector(to_unsigned( 116,8)),
			13914 => std_logic_vector(to_unsigned( 176,8)),
			13915 => std_logic_vector(to_unsigned( 114,8)),
			13916 => std_logic_vector(to_unsigned( 251,8)),
			13917 => std_logic_vector(to_unsigned( 166,8)),
			13918 => std_logic_vector(to_unsigned( 53,8)),
			13919 => std_logic_vector(to_unsigned( 22,8)),
			13920 => std_logic_vector(to_unsigned( 80,8)),
			13921 => std_logic_vector(to_unsigned( 95,8)),
			13922 => std_logic_vector(to_unsigned( 219,8)),
			13923 => std_logic_vector(to_unsigned( 108,8)),
			13924 => std_logic_vector(to_unsigned( 15,8)),
			13925 => std_logic_vector(to_unsigned( 77,8)),
			13926 => std_logic_vector(to_unsigned( 156,8)),
			13927 => std_logic_vector(to_unsigned( 169,8)),
			13928 => std_logic_vector(to_unsigned( 27,8)),
			13929 => std_logic_vector(to_unsigned( 164,8)),
			13930 => std_logic_vector(to_unsigned( 118,8)),
			13931 => std_logic_vector(to_unsigned( 33,8)),
			13932 => std_logic_vector(to_unsigned( 159,8)),
			13933 => std_logic_vector(to_unsigned( 167,8)),
			13934 => std_logic_vector(to_unsigned( 8,8)),
			13935 => std_logic_vector(to_unsigned( 124,8)),
			13936 => std_logic_vector(to_unsigned( 106,8)),
			13937 => std_logic_vector(to_unsigned( 174,8)),
			13938 => std_logic_vector(to_unsigned( 173,8)),
			13939 => std_logic_vector(to_unsigned( 250,8)),
			13940 => std_logic_vector(to_unsigned( 186,8)),
			13941 => std_logic_vector(to_unsigned( 194,8)),
			13942 => std_logic_vector(to_unsigned( 74,8)),
			13943 => std_logic_vector(to_unsigned( 40,8)),
			13944 => std_logic_vector(to_unsigned( 70,8)),
			13945 => std_logic_vector(to_unsigned( 15,8)),
			13946 => std_logic_vector(to_unsigned( 117,8)),
			13947 => std_logic_vector(to_unsigned( 122,8)),
			13948 => std_logic_vector(to_unsigned( 170,8)),
			13949 => std_logic_vector(to_unsigned( 175,8)),
			13950 => std_logic_vector(to_unsigned( 46,8)),
			13951 => std_logic_vector(to_unsigned( 195,8)),
			13952 => std_logic_vector(to_unsigned( 53,8)),
			13953 => std_logic_vector(to_unsigned( 225,8)),
			13954 => std_logic_vector(to_unsigned( 36,8)),
			13955 => std_logic_vector(to_unsigned( 164,8)),
			13956 => std_logic_vector(to_unsigned( 227,8)),
			13957 => std_logic_vector(to_unsigned( 239,8)),
			13958 => std_logic_vector(to_unsigned( 150,8)),
			13959 => std_logic_vector(to_unsigned( 242,8)),
			13960 => std_logic_vector(to_unsigned( 85,8)),
			13961 => std_logic_vector(to_unsigned( 16,8)),
			13962 => std_logic_vector(to_unsigned( 68,8)),
			13963 => std_logic_vector(to_unsigned( 3,8)),
			13964 => std_logic_vector(to_unsigned( 59,8)),
			13965 => std_logic_vector(to_unsigned( 248,8)),
			13966 => std_logic_vector(to_unsigned( 227,8)),
			13967 => std_logic_vector(to_unsigned( 226,8)),
			13968 => std_logic_vector(to_unsigned( 213,8)),
			13969 => std_logic_vector(to_unsigned( 117,8)),
			13970 => std_logic_vector(to_unsigned( 151,8)),
			13971 => std_logic_vector(to_unsigned( 18,8)),
			13972 => std_logic_vector(to_unsigned( 138,8)),
			13973 => std_logic_vector(to_unsigned( 114,8)),
			13974 => std_logic_vector(to_unsigned( 143,8)),
			13975 => std_logic_vector(to_unsigned( 97,8)),
			13976 => std_logic_vector(to_unsigned( 73,8)),
			13977 => std_logic_vector(to_unsigned( 242,8)),
			13978 => std_logic_vector(to_unsigned( 158,8)),
			13979 => std_logic_vector(to_unsigned( 10,8)),
			13980 => std_logic_vector(to_unsigned( 73,8)),
			13981 => std_logic_vector(to_unsigned( 55,8)),
			13982 => std_logic_vector(to_unsigned( 73,8)),
			13983 => std_logic_vector(to_unsigned( 142,8)),
			13984 => std_logic_vector(to_unsigned( 137,8)),
			13985 => std_logic_vector(to_unsigned( 253,8)),
			13986 => std_logic_vector(to_unsigned( 13,8)),
			13987 => std_logic_vector(to_unsigned( 127,8)),
			13988 => std_logic_vector(to_unsigned( 55,8)),
			13989 => std_logic_vector(to_unsigned( 58,8)),
			13990 => std_logic_vector(to_unsigned( 77,8)),
			13991 => std_logic_vector(to_unsigned( 4,8)),
			13992 => std_logic_vector(to_unsigned( 124,8)),
			13993 => std_logic_vector(to_unsigned( 83,8)),
			13994 => std_logic_vector(to_unsigned( 184,8)),
			13995 => std_logic_vector(to_unsigned( 123,8)),
			13996 => std_logic_vector(to_unsigned( 106,8)),
			13997 => std_logic_vector(to_unsigned( 160,8)),
			13998 => std_logic_vector(to_unsigned( 132,8)),
			13999 => std_logic_vector(to_unsigned( 68,8)),
			14000 => std_logic_vector(to_unsigned( 38,8)),
			14001 => std_logic_vector(to_unsigned( 57,8)),
			14002 => std_logic_vector(to_unsigned( 109,8)),
			14003 => std_logic_vector(to_unsigned( 141,8)),
			14004 => std_logic_vector(to_unsigned( 221,8)),
			14005 => std_logic_vector(to_unsigned( 198,8)),
			14006 => std_logic_vector(to_unsigned( 39,8)),
			14007 => std_logic_vector(to_unsigned( 182,8)),
			14008 => std_logic_vector(to_unsigned( 102,8)),
			14009 => std_logic_vector(to_unsigned( 225,8)),
			14010 => std_logic_vector(to_unsigned( 228,8)),
			14011 => std_logic_vector(to_unsigned( 10,8)),
			14012 => std_logic_vector(to_unsigned( 9,8)),
			14013 => std_logic_vector(to_unsigned( 210,8)),
			14014 => std_logic_vector(to_unsigned( 25,8)),
			14015 => std_logic_vector(to_unsigned( 133,8)),
			14016 => std_logic_vector(to_unsigned( 207,8)),
			14017 => std_logic_vector(to_unsigned( 139,8)),
			14018 => std_logic_vector(to_unsigned( 75,8)),
			14019 => std_logic_vector(to_unsigned( 164,8)),
			14020 => std_logic_vector(to_unsigned( 83,8)),
			14021 => std_logic_vector(to_unsigned( 12,8)),
			14022 => std_logic_vector(to_unsigned( 227,8)),
			14023 => std_logic_vector(to_unsigned( 234,8)),
			14024 => std_logic_vector(to_unsigned( 70,8)),
			14025 => std_logic_vector(to_unsigned( 198,8)),
			14026 => std_logic_vector(to_unsigned( 182,8)),
			14027 => std_logic_vector(to_unsigned( 29,8)),
			14028 => std_logic_vector(to_unsigned( 197,8)),
			14029 => std_logic_vector(to_unsigned( 105,8)),
			14030 => std_logic_vector(to_unsigned( 74,8)),
			14031 => std_logic_vector(to_unsigned( 73,8)),
			14032 => std_logic_vector(to_unsigned( 59,8)),
			14033 => std_logic_vector(to_unsigned( 0,8)),
			14034 => std_logic_vector(to_unsigned( 169,8)),
			14035 => std_logic_vector(to_unsigned( 94,8)),
			14036 => std_logic_vector(to_unsigned( 139,8)),
			14037 => std_logic_vector(to_unsigned( 244,8)),
			14038 => std_logic_vector(to_unsigned( 135,8)),
			14039 => std_logic_vector(to_unsigned( 185,8)),
			14040 => std_logic_vector(to_unsigned( 88,8)),
			14041 => std_logic_vector(to_unsigned( 240,8)),
			14042 => std_logic_vector(to_unsigned( 249,8)),
			14043 => std_logic_vector(to_unsigned( 253,8)),
			14044 => std_logic_vector(to_unsigned( 156,8)),
			14045 => std_logic_vector(to_unsigned( 71,8)),
			14046 => std_logic_vector(to_unsigned( 212,8)),
			14047 => std_logic_vector(to_unsigned( 72,8)),
			14048 => std_logic_vector(to_unsigned( 144,8)),
			14049 => std_logic_vector(to_unsigned( 30,8)),
			14050 => std_logic_vector(to_unsigned( 87,8)),
			14051 => std_logic_vector(to_unsigned( 109,8)),
			14052 => std_logic_vector(to_unsigned( 196,8)),
			14053 => std_logic_vector(to_unsigned( 88,8)),
			14054 => std_logic_vector(to_unsigned( 100,8)),
			14055 => std_logic_vector(to_unsigned( 46,8)),
			14056 => std_logic_vector(to_unsigned( 120,8)),
			14057 => std_logic_vector(to_unsigned( 106,8)),
			14058 => std_logic_vector(to_unsigned( 244,8)),
			14059 => std_logic_vector(to_unsigned( 44,8)),
			14060 => std_logic_vector(to_unsigned( 11,8)),
			14061 => std_logic_vector(to_unsigned( 158,8)),
			14062 => std_logic_vector(to_unsigned( 52,8)),
			14063 => std_logic_vector(to_unsigned( 56,8)),
			14064 => std_logic_vector(to_unsigned( 174,8)),
			14065 => std_logic_vector(to_unsigned( 0,8)),
			14066 => std_logic_vector(to_unsigned( 110,8)),
			14067 => std_logic_vector(to_unsigned( 126,8)),
			14068 => std_logic_vector(to_unsigned( 210,8)),
			14069 => std_logic_vector(to_unsigned( 45,8)),
			14070 => std_logic_vector(to_unsigned( 159,8)),
			14071 => std_logic_vector(to_unsigned( 245,8)),
			14072 => std_logic_vector(to_unsigned( 198,8)),
			14073 => std_logic_vector(to_unsigned( 74,8)),
			14074 => std_logic_vector(to_unsigned( 207,8)),
			14075 => std_logic_vector(to_unsigned( 26,8)),
			14076 => std_logic_vector(to_unsigned( 54,8)),
			14077 => std_logic_vector(to_unsigned( 212,8)),
			14078 => std_logic_vector(to_unsigned( 89,8)),
			14079 => std_logic_vector(to_unsigned( 108,8)),
			14080 => std_logic_vector(to_unsigned( 182,8)),
			14081 => std_logic_vector(to_unsigned( 229,8)),
			14082 => std_logic_vector(to_unsigned( 235,8)),
			14083 => std_logic_vector(to_unsigned( 224,8)),
			14084 => std_logic_vector(to_unsigned( 172,8)),
			14085 => std_logic_vector(to_unsigned( 137,8)),
			14086 => std_logic_vector(to_unsigned( 230,8)),
			14087 => std_logic_vector(to_unsigned( 154,8)),
			14088 => std_logic_vector(to_unsigned( 151,8)),
			14089 => std_logic_vector(to_unsigned( 119,8)),
			14090 => std_logic_vector(to_unsigned( 8,8)),
			14091 => std_logic_vector(to_unsigned( 19,8)),
			14092 => std_logic_vector(to_unsigned( 160,8)),
			14093 => std_logic_vector(to_unsigned( 26,8)),
			14094 => std_logic_vector(to_unsigned( 5,8)),
			14095 => std_logic_vector(to_unsigned( 202,8)),
			14096 => std_logic_vector(to_unsigned( 72,8)),
			14097 => std_logic_vector(to_unsigned( 31,8)),
			14098 => std_logic_vector(to_unsigned( 142,8)),
			14099 => std_logic_vector(to_unsigned( 20,8)),
			14100 => std_logic_vector(to_unsigned( 111,8)),
			14101 => std_logic_vector(to_unsigned( 188,8)),
			14102 => std_logic_vector(to_unsigned( 57,8)),
			14103 => std_logic_vector(to_unsigned( 134,8)),
			14104 => std_logic_vector(to_unsigned( 81,8)),
			14105 => std_logic_vector(to_unsigned( 40,8)),
			14106 => std_logic_vector(to_unsigned( 33,8)),
			14107 => std_logic_vector(to_unsigned( 42,8)),
			14108 => std_logic_vector(to_unsigned( 68,8)),
			14109 => std_logic_vector(to_unsigned( 26,8)),
			14110 => std_logic_vector(to_unsigned( 200,8)),
			14111 => std_logic_vector(to_unsigned( 81,8)),
			14112 => std_logic_vector(to_unsigned( 105,8)),
			14113 => std_logic_vector(to_unsigned( 23,8)),
			14114 => std_logic_vector(to_unsigned( 254,8)),
			14115 => std_logic_vector(to_unsigned( 141,8)),
			14116 => std_logic_vector(to_unsigned( 21,8)),
			14117 => std_logic_vector(to_unsigned( 195,8)),
			14118 => std_logic_vector(to_unsigned( 174,8)),
			14119 => std_logic_vector(to_unsigned( 249,8)),
			14120 => std_logic_vector(to_unsigned( 55,8)),
			14121 => std_logic_vector(to_unsigned( 112,8)),
			14122 => std_logic_vector(to_unsigned( 26,8)),
			14123 => std_logic_vector(to_unsigned( 79,8)),
			14124 => std_logic_vector(to_unsigned( 119,8)),
			14125 => std_logic_vector(to_unsigned( 27,8)),
			14126 => std_logic_vector(to_unsigned( 126,8)),
			14127 => std_logic_vector(to_unsigned( 51,8)),
			14128 => std_logic_vector(to_unsigned( 212,8)),
			14129 => std_logic_vector(to_unsigned( 147,8)),
			14130 => std_logic_vector(to_unsigned( 143,8)),
			14131 => std_logic_vector(to_unsigned( 151,8)),
			14132 => std_logic_vector(to_unsigned( 73,8)),
			14133 => std_logic_vector(to_unsigned( 23,8)),
			14134 => std_logic_vector(to_unsigned( 250,8)),
			14135 => std_logic_vector(to_unsigned( 202,8)),
			14136 => std_logic_vector(to_unsigned( 73,8)),
			14137 => std_logic_vector(to_unsigned( 127,8)),
			14138 => std_logic_vector(to_unsigned( 117,8)),
			14139 => std_logic_vector(to_unsigned( 67,8)),
			14140 => std_logic_vector(to_unsigned( 198,8)),
			14141 => std_logic_vector(to_unsigned( 214,8)),
			14142 => std_logic_vector(to_unsigned( 134,8)),
			14143 => std_logic_vector(to_unsigned( 19,8)),
			14144 => std_logic_vector(to_unsigned( 123,8)),
			14145 => std_logic_vector(to_unsigned( 59,8)),
			14146 => std_logic_vector(to_unsigned( 21,8)),
			14147 => std_logic_vector(to_unsigned( 239,8)),
			14148 => std_logic_vector(to_unsigned( 16,8)),
			14149 => std_logic_vector(to_unsigned( 126,8)),
			14150 => std_logic_vector(to_unsigned( 63,8)),
			14151 => std_logic_vector(to_unsigned( 88,8)),
			14152 => std_logic_vector(to_unsigned( 133,8)),
			14153 => std_logic_vector(to_unsigned( 28,8)),
			14154 => std_logic_vector(to_unsigned( 235,8)),
			14155 => std_logic_vector(to_unsigned( 44,8)),
			14156 => std_logic_vector(to_unsigned( 172,8)),
			14157 => std_logic_vector(to_unsigned( 101,8)),
			14158 => std_logic_vector(to_unsigned( 136,8)),
			14159 => std_logic_vector(to_unsigned( 158,8)),
			14160 => std_logic_vector(to_unsigned( 38,8)),
			14161 => std_logic_vector(to_unsigned( 97,8)),
			14162 => std_logic_vector(to_unsigned( 174,8)),
			14163 => std_logic_vector(to_unsigned( 46,8)),
			14164 => std_logic_vector(to_unsigned( 97,8)),
			14165 => std_logic_vector(to_unsigned( 132,8)),
			14166 => std_logic_vector(to_unsigned( 228,8)),
			14167 => std_logic_vector(to_unsigned( 213,8)),
			14168 => std_logic_vector(to_unsigned( 170,8)),
			14169 => std_logic_vector(to_unsigned( 37,8)),
			14170 => std_logic_vector(to_unsigned( 245,8)),
			14171 => std_logic_vector(to_unsigned( 5,8)),
			14172 => std_logic_vector(to_unsigned( 9,8)),
			14173 => std_logic_vector(to_unsigned( 164,8)),
			14174 => std_logic_vector(to_unsigned( 39,8)),
			14175 => std_logic_vector(to_unsigned( 117,8)),
			14176 => std_logic_vector(to_unsigned( 55,8)),
			14177 => std_logic_vector(to_unsigned( 200,8)),
			14178 => std_logic_vector(to_unsigned( 180,8)),
			14179 => std_logic_vector(to_unsigned( 126,8)),
			14180 => std_logic_vector(to_unsigned( 193,8)),
			14181 => std_logic_vector(to_unsigned( 70,8)),
			14182 => std_logic_vector(to_unsigned( 235,8)),
			14183 => std_logic_vector(to_unsigned( 68,8)),
			14184 => std_logic_vector(to_unsigned( 70,8)),
			14185 => std_logic_vector(to_unsigned( 16,8)),
			14186 => std_logic_vector(to_unsigned( 126,8)),
			14187 => std_logic_vector(to_unsigned( 205,8)),
			14188 => std_logic_vector(to_unsigned( 53,8)),
			14189 => std_logic_vector(to_unsigned( 234,8)),
			14190 => std_logic_vector(to_unsigned( 161,8)),
			14191 => std_logic_vector(to_unsigned( 244,8)),
			14192 => std_logic_vector(to_unsigned( 209,8)),
			14193 => std_logic_vector(to_unsigned( 111,8)),
			14194 => std_logic_vector(to_unsigned( 15,8)),
			14195 => std_logic_vector(to_unsigned( 51,8)),
			14196 => std_logic_vector(to_unsigned( 33,8)),
			14197 => std_logic_vector(to_unsigned( 120,8)),
			14198 => std_logic_vector(to_unsigned( 54,8)),
			14199 => std_logic_vector(to_unsigned( 40,8)),
			14200 => std_logic_vector(to_unsigned( 95,8)),
			14201 => std_logic_vector(to_unsigned( 226,8)),
			14202 => std_logic_vector(to_unsigned( 156,8)),
			14203 => std_logic_vector(to_unsigned( 115,8)),
			14204 => std_logic_vector(to_unsigned( 25,8)),
			14205 => std_logic_vector(to_unsigned( 235,8)),
			14206 => std_logic_vector(to_unsigned( 143,8)),
			14207 => std_logic_vector(to_unsigned( 225,8)),
			14208 => std_logic_vector(to_unsigned( 92,8)),
			14209 => std_logic_vector(to_unsigned( 25,8)),
			14210 => std_logic_vector(to_unsigned( 198,8)),
			14211 => std_logic_vector(to_unsigned( 146,8)),
			14212 => std_logic_vector(to_unsigned( 19,8)),
			14213 => std_logic_vector(to_unsigned( 220,8)),
			14214 => std_logic_vector(to_unsigned( 89,8)),
			14215 => std_logic_vector(to_unsigned( 221,8)),
			14216 => std_logic_vector(to_unsigned( 245,8)),
			14217 => std_logic_vector(to_unsigned( 129,8)),
			14218 => std_logic_vector(to_unsigned( 190,8)),
			14219 => std_logic_vector(to_unsigned( 11,8)),
			14220 => std_logic_vector(to_unsigned( 210,8)),
			14221 => std_logic_vector(to_unsigned( 22,8)),
			14222 => std_logic_vector(to_unsigned( 218,8)),
			14223 => std_logic_vector(to_unsigned( 231,8)),
			14224 => std_logic_vector(to_unsigned( 129,8)),
			14225 => std_logic_vector(to_unsigned( 161,8)),
			14226 => std_logic_vector(to_unsigned( 227,8)),
			14227 => std_logic_vector(to_unsigned( 55,8)),
			14228 => std_logic_vector(to_unsigned( 153,8)),
			14229 => std_logic_vector(to_unsigned( 88,8)),
			14230 => std_logic_vector(to_unsigned( 69,8)),
			14231 => std_logic_vector(to_unsigned( 55,8)),
			14232 => std_logic_vector(to_unsigned( 185,8)),
			14233 => std_logic_vector(to_unsigned( 46,8)),
			14234 => std_logic_vector(to_unsigned( 134,8)),
			14235 => std_logic_vector(to_unsigned( 114,8)),
			14236 => std_logic_vector(to_unsigned( 29,8)),
			14237 => std_logic_vector(to_unsigned( 76,8)),
			14238 => std_logic_vector(to_unsigned( 20,8)),
			14239 => std_logic_vector(to_unsigned( 155,8)),
			14240 => std_logic_vector(to_unsigned( 49,8)),
			14241 => std_logic_vector(to_unsigned( 207,8)),
			14242 => std_logic_vector(to_unsigned( 166,8)),
			14243 => std_logic_vector(to_unsigned( 120,8)),
			14244 => std_logic_vector(to_unsigned( 3,8)),
			14245 => std_logic_vector(to_unsigned( 235,8)),
			14246 => std_logic_vector(to_unsigned( 194,8)),
			14247 => std_logic_vector(to_unsigned( 92,8)),
			14248 => std_logic_vector(to_unsigned( 197,8)),
			14249 => std_logic_vector(to_unsigned( 110,8)),
			14250 => std_logic_vector(to_unsigned( 114,8)),
			14251 => std_logic_vector(to_unsigned( 57,8)),
			14252 => std_logic_vector(to_unsigned( 171,8)),
			14253 => std_logic_vector(to_unsigned( 223,8)),
			14254 => std_logic_vector(to_unsigned( 204,8)),
			14255 => std_logic_vector(to_unsigned( 51,8)),
			14256 => std_logic_vector(to_unsigned( 114,8)),
			14257 => std_logic_vector(to_unsigned( 208,8)),
			14258 => std_logic_vector(to_unsigned( 141,8)),
			14259 => std_logic_vector(to_unsigned( 220,8)),
			14260 => std_logic_vector(to_unsigned( 238,8)),
			14261 => std_logic_vector(to_unsigned( 106,8)),
			14262 => std_logic_vector(to_unsigned( 4,8)),
			14263 => std_logic_vector(to_unsigned( 61,8)),
			14264 => std_logic_vector(to_unsigned( 166,8)),
			14265 => std_logic_vector(to_unsigned( 214,8)),
			14266 => std_logic_vector(to_unsigned( 207,8)),
			14267 => std_logic_vector(to_unsigned( 254,8)),
			14268 => std_logic_vector(to_unsigned( 27,8)),
			14269 => std_logic_vector(to_unsigned( 186,8)),
			14270 => std_logic_vector(to_unsigned( 74,8)),
			14271 => std_logic_vector(to_unsigned( 24,8)),
			14272 => std_logic_vector(to_unsigned( 170,8)),
			14273 => std_logic_vector(to_unsigned( 67,8)),
			14274 => std_logic_vector(to_unsigned( 85,8)),
			14275 => std_logic_vector(to_unsigned( 204,8)),
			14276 => std_logic_vector(to_unsigned( 69,8)),
			14277 => std_logic_vector(to_unsigned( 51,8)),
			14278 => std_logic_vector(to_unsigned( 123,8)),
			14279 => std_logic_vector(to_unsigned( 82,8)),
			14280 => std_logic_vector(to_unsigned( 219,8)),
			14281 => std_logic_vector(to_unsigned( 237,8)),
			14282 => std_logic_vector(to_unsigned( 119,8)),
			14283 => std_logic_vector(to_unsigned( 37,8)),
			14284 => std_logic_vector(to_unsigned( 17,8)),
			14285 => std_logic_vector(to_unsigned( 87,8)),
			14286 => std_logic_vector(to_unsigned( 108,8)),
			14287 => std_logic_vector(to_unsigned( 131,8)),
			14288 => std_logic_vector(to_unsigned( 159,8)),
			14289 => std_logic_vector(to_unsigned( 83,8)),
			14290 => std_logic_vector(to_unsigned( 181,8)),
			14291 => std_logic_vector(to_unsigned( 216,8)),
			14292 => std_logic_vector(to_unsigned( 38,8)),
			14293 => std_logic_vector(to_unsigned( 218,8)),
			14294 => std_logic_vector(to_unsigned( 49,8)),
			14295 => std_logic_vector(to_unsigned( 120,8)),
			14296 => std_logic_vector(to_unsigned( 25,8)),
			14297 => std_logic_vector(to_unsigned( 174,8)),
			14298 => std_logic_vector(to_unsigned( 147,8)),
			14299 => std_logic_vector(to_unsigned( 195,8)),
			14300 => std_logic_vector(to_unsigned( 172,8)),
			14301 => std_logic_vector(to_unsigned( 76,8)),
			14302 => std_logic_vector(to_unsigned( 33,8)),
			14303 => std_logic_vector(to_unsigned( 72,8)),
			14304 => std_logic_vector(to_unsigned( 128,8)),
			14305 => std_logic_vector(to_unsigned( 86,8)),
			14306 => std_logic_vector(to_unsigned( 236,8)),
			14307 => std_logic_vector(to_unsigned( 254,8)),
			14308 => std_logic_vector(to_unsigned( 183,8)),
			14309 => std_logic_vector(to_unsigned( 239,8)),
			14310 => std_logic_vector(to_unsigned( 172,8)),
			14311 => std_logic_vector(to_unsigned( 92,8)),
			14312 => std_logic_vector(to_unsigned( 3,8)),
			14313 => std_logic_vector(to_unsigned( 7,8)),
			14314 => std_logic_vector(to_unsigned( 165,8)),
			14315 => std_logic_vector(to_unsigned( 174,8)),
			14316 => std_logic_vector(to_unsigned( 166,8)),
			14317 => std_logic_vector(to_unsigned( 184,8)),
			14318 => std_logic_vector(to_unsigned( 147,8)),
			14319 => std_logic_vector(to_unsigned( 181,8)),
			14320 => std_logic_vector(to_unsigned( 30,8)),
			14321 => std_logic_vector(to_unsigned( 199,8)),
			14322 => std_logic_vector(to_unsigned( 101,8)),
			14323 => std_logic_vector(to_unsigned( 200,8)),
			14324 => std_logic_vector(to_unsigned( 129,8)),
			14325 => std_logic_vector(to_unsigned( 131,8)),
			14326 => std_logic_vector(to_unsigned( 81,8)),
			14327 => std_logic_vector(to_unsigned( 230,8)),
			14328 => std_logic_vector(to_unsigned( 53,8)),
			14329 => std_logic_vector(to_unsigned( 114,8)),
			14330 => std_logic_vector(to_unsigned( 2,8)),
			14331 => std_logic_vector(to_unsigned( 232,8)),
			14332 => std_logic_vector(to_unsigned( 212,8)),
			14333 => std_logic_vector(to_unsigned( 96,8)),
			14334 => std_logic_vector(to_unsigned( 196,8)),
			14335 => std_logic_vector(to_unsigned( 66,8)),
			14336 => std_logic_vector(to_unsigned( 18,8)),
			14337 => std_logic_vector(to_unsigned( 84,8)),
			14338 => std_logic_vector(to_unsigned( 103,8)),
			14339 => std_logic_vector(to_unsigned( 4,8)),
			14340 => std_logic_vector(to_unsigned( 78,8)),
			14341 => std_logic_vector(to_unsigned( 119,8)),
			14342 => std_logic_vector(to_unsigned( 23,8)),
			14343 => std_logic_vector(to_unsigned( 119,8)),
			14344 => std_logic_vector(to_unsigned( 71,8)),
			14345 => std_logic_vector(to_unsigned( 125,8)),
			14346 => std_logic_vector(to_unsigned( 113,8)),
			14347 => std_logic_vector(to_unsigned( 13,8)),
			14348 => std_logic_vector(to_unsigned( 54,8)),
			14349 => std_logic_vector(to_unsigned( 135,8)),
			14350 => std_logic_vector(to_unsigned( 143,8)),
			14351 => std_logic_vector(to_unsigned( 250,8)),
			14352 => std_logic_vector(to_unsigned( 86,8)),
			14353 => std_logic_vector(to_unsigned( 169,8)),
			14354 => std_logic_vector(to_unsigned( 7,8)),
			14355 => std_logic_vector(to_unsigned( 117,8)),
			14356 => std_logic_vector(to_unsigned( 110,8)),
			14357 => std_logic_vector(to_unsigned( 58,8)),
			14358 => std_logic_vector(to_unsigned( 81,8)),
			14359 => std_logic_vector(to_unsigned( 22,8)),
			14360 => std_logic_vector(to_unsigned( 247,8)),
			14361 => std_logic_vector(to_unsigned( 112,8)),
			14362 => std_logic_vector(to_unsigned( 78,8)),
			14363 => std_logic_vector(to_unsigned( 4,8)),
			14364 => std_logic_vector(to_unsigned( 18,8)),
			14365 => std_logic_vector(to_unsigned( 32,8)),
			14366 => std_logic_vector(to_unsigned( 17,8)),
			14367 => std_logic_vector(to_unsigned( 218,8)),
			14368 => std_logic_vector(to_unsigned( 155,8)),
			14369 => std_logic_vector(to_unsigned( 212,8)),
			14370 => std_logic_vector(to_unsigned( 90,8)),
			14371 => std_logic_vector(to_unsigned( 97,8)),
			14372 => std_logic_vector(to_unsigned( 20,8)),
			14373 => std_logic_vector(to_unsigned( 111,8)),
			14374 => std_logic_vector(to_unsigned( 88,8)),
			14375 => std_logic_vector(to_unsigned( 210,8)),
			14376 => std_logic_vector(to_unsigned( 100,8)),
			14377 => std_logic_vector(to_unsigned( 17,8)),
			14378 => std_logic_vector(to_unsigned( 140,8)),
			14379 => std_logic_vector(to_unsigned( 16,8)),
			14380 => std_logic_vector(to_unsigned( 233,8)),
			14381 => std_logic_vector(to_unsigned( 215,8)),
			14382 => std_logic_vector(to_unsigned( 126,8)),
			14383 => std_logic_vector(to_unsigned( 179,8)),
			14384 => std_logic_vector(to_unsigned( 163,8)),
			14385 => std_logic_vector(to_unsigned( 222,8)),
			14386 => std_logic_vector(to_unsigned( 144,8)),
			14387 => std_logic_vector(to_unsigned( 83,8)),
			14388 => std_logic_vector(to_unsigned( 173,8)),
			14389 => std_logic_vector(to_unsigned( 218,8)),
			14390 => std_logic_vector(to_unsigned( 167,8)),
			14391 => std_logic_vector(to_unsigned( 109,8)),
			14392 => std_logic_vector(to_unsigned( 140,8)),
			14393 => std_logic_vector(to_unsigned( 11,8)),
			14394 => std_logic_vector(to_unsigned( 155,8)),
			14395 => std_logic_vector(to_unsigned( 59,8)),
			14396 => std_logic_vector(to_unsigned( 75,8)),
			14397 => std_logic_vector(to_unsigned( 221,8)),
			14398 => std_logic_vector(to_unsigned( 213,8)),
			14399 => std_logic_vector(to_unsigned( 53,8)),
			14400 => std_logic_vector(to_unsigned( 115,8)),
			14401 => std_logic_vector(to_unsigned( 26,8)),
			14402 => std_logic_vector(to_unsigned( 156,8)),
			14403 => std_logic_vector(to_unsigned( 8,8)),
			14404 => std_logic_vector(to_unsigned( 2,8)),
			14405 => std_logic_vector(to_unsigned( 229,8)),
			14406 => std_logic_vector(to_unsigned( 99,8)),
			14407 => std_logic_vector(to_unsigned( 214,8)),
			14408 => std_logic_vector(to_unsigned( 219,8)),
			14409 => std_logic_vector(to_unsigned( 8,8)),
			14410 => std_logic_vector(to_unsigned( 113,8)),
			14411 => std_logic_vector(to_unsigned( 40,8)),
			14412 => std_logic_vector(to_unsigned( 48,8)),
			14413 => std_logic_vector(to_unsigned( 249,8)),
			14414 => std_logic_vector(to_unsigned( 55,8)),
			14415 => std_logic_vector(to_unsigned( 47,8)),
			14416 => std_logic_vector(to_unsigned( 57,8)),
			14417 => std_logic_vector(to_unsigned( 143,8)),
			14418 => std_logic_vector(to_unsigned( 137,8)),
			14419 => std_logic_vector(to_unsigned( 181,8)),
			14420 => std_logic_vector(to_unsigned( 172,8)),
			14421 => std_logic_vector(to_unsigned( 139,8)),
			14422 => std_logic_vector(to_unsigned( 58,8)),
			14423 => std_logic_vector(to_unsigned( 100,8)),
			14424 => std_logic_vector(to_unsigned( 39,8)),
			14425 => std_logic_vector(to_unsigned( 255,8)),
			14426 => std_logic_vector(to_unsigned( 170,8)),
			14427 => std_logic_vector(to_unsigned( 86,8)),
			14428 => std_logic_vector(to_unsigned( 252,8)),
			14429 => std_logic_vector(to_unsigned( 251,8)),
			14430 => std_logic_vector(to_unsigned( 109,8)),
			14431 => std_logic_vector(to_unsigned( 51,8)),
			14432 => std_logic_vector(to_unsigned( 18,8)),
			14433 => std_logic_vector(to_unsigned( 112,8)),
			14434 => std_logic_vector(to_unsigned( 128,8)),
			14435 => std_logic_vector(to_unsigned( 218,8)),
			14436 => std_logic_vector(to_unsigned( 252,8)),
			14437 => std_logic_vector(to_unsigned( 183,8)),
			14438 => std_logic_vector(to_unsigned( 81,8)),
			14439 => std_logic_vector(to_unsigned( 142,8)),
			14440 => std_logic_vector(to_unsigned( 106,8)),
			14441 => std_logic_vector(to_unsigned( 63,8)),
			14442 => std_logic_vector(to_unsigned( 192,8)),
			14443 => std_logic_vector(to_unsigned( 24,8)),
			14444 => std_logic_vector(to_unsigned( 5,8)),
			14445 => std_logic_vector(to_unsigned( 24,8)),
			14446 => std_logic_vector(to_unsigned( 92,8)),
			14447 => std_logic_vector(to_unsigned( 105,8)),
			14448 => std_logic_vector(to_unsigned( 111,8)),
			14449 => std_logic_vector(to_unsigned( 253,8)),
			14450 => std_logic_vector(to_unsigned( 69,8)),
			14451 => std_logic_vector(to_unsigned( 217,8)),
			14452 => std_logic_vector(to_unsigned( 174,8)),
			14453 => std_logic_vector(to_unsigned( 135,8)),
			14454 => std_logic_vector(to_unsigned( 204,8)),
			14455 => std_logic_vector(to_unsigned( 243,8)),
			14456 => std_logic_vector(to_unsigned( 140,8)),
			14457 => std_logic_vector(to_unsigned( 174,8)),
			14458 => std_logic_vector(to_unsigned( 249,8)),
			14459 => std_logic_vector(to_unsigned( 246,8)),
			14460 => std_logic_vector(to_unsigned( 29,8)),
			14461 => std_logic_vector(to_unsigned( 79,8)),
			14462 => std_logic_vector(to_unsigned( 14,8)),
			14463 => std_logic_vector(to_unsigned( 51,8)),
			14464 => std_logic_vector(to_unsigned( 77,8)),
			14465 => std_logic_vector(to_unsigned( 86,8)),
			14466 => std_logic_vector(to_unsigned( 252,8)),
			14467 => std_logic_vector(to_unsigned( 243,8)),
			14468 => std_logic_vector(to_unsigned( 97,8)),
			14469 => std_logic_vector(to_unsigned( 2,8)),
			14470 => std_logic_vector(to_unsigned( 82,8)),
			14471 => std_logic_vector(to_unsigned( 181,8)),
			14472 => std_logic_vector(to_unsigned( 99,8)),
			14473 => std_logic_vector(to_unsigned( 99,8)),
			14474 => std_logic_vector(to_unsigned( 72,8)),
			14475 => std_logic_vector(to_unsigned( 29,8)),
			14476 => std_logic_vector(to_unsigned( 234,8)),
			14477 => std_logic_vector(to_unsigned( 147,8)),
			14478 => std_logic_vector(to_unsigned( 133,8)),
			14479 => std_logic_vector(to_unsigned( 191,8)),
			14480 => std_logic_vector(to_unsigned( 52,8)),
			14481 => std_logic_vector(to_unsigned( 139,8)),
			14482 => std_logic_vector(to_unsigned( 237,8)),
			14483 => std_logic_vector(to_unsigned( 190,8)),
			14484 => std_logic_vector(to_unsigned( 183,8)),
			14485 => std_logic_vector(to_unsigned( 197,8)),
			14486 => std_logic_vector(to_unsigned( 42,8)),
			14487 => std_logic_vector(to_unsigned( 55,8)),
			14488 => std_logic_vector(to_unsigned( 160,8)),
			14489 => std_logic_vector(to_unsigned( 114,8)),
			14490 => std_logic_vector(to_unsigned( 154,8)),
			14491 => std_logic_vector(to_unsigned( 179,8)),
			14492 => std_logic_vector(to_unsigned( 228,8)),
			14493 => std_logic_vector(to_unsigned( 156,8)),
			14494 => std_logic_vector(to_unsigned( 116,8)),
			14495 => std_logic_vector(to_unsigned( 58,8)),
			14496 => std_logic_vector(to_unsigned( 238,8)),
			14497 => std_logic_vector(to_unsigned( 253,8)),
			14498 => std_logic_vector(to_unsigned( 179,8)),
			14499 => std_logic_vector(to_unsigned( 241,8)),
			14500 => std_logic_vector(to_unsigned( 51,8)),
			14501 => std_logic_vector(to_unsigned( 246,8)),
			14502 => std_logic_vector(to_unsigned( 123,8)),
			14503 => std_logic_vector(to_unsigned( 23,8)),
			14504 => std_logic_vector(to_unsigned( 238,8)),
			14505 => std_logic_vector(to_unsigned( 162,8)),
			14506 => std_logic_vector(to_unsigned( 29,8)),
			14507 => std_logic_vector(to_unsigned( 132,8)),
			14508 => std_logic_vector(to_unsigned( 101,8)),
			14509 => std_logic_vector(to_unsigned( 199,8)),
			14510 => std_logic_vector(to_unsigned( 238,8)),
			14511 => std_logic_vector(to_unsigned( 210,8)),
			14512 => std_logic_vector(to_unsigned( 198,8)),
			14513 => std_logic_vector(to_unsigned( 169,8)),
			14514 => std_logic_vector(to_unsigned( 239,8)),
			14515 => std_logic_vector(to_unsigned( 22,8)),
			14516 => std_logic_vector(to_unsigned( 223,8)),
			14517 => std_logic_vector(to_unsigned( 61,8)),
			14518 => std_logic_vector(to_unsigned( 72,8)),
			14519 => std_logic_vector(to_unsigned( 80,8)),
			14520 => std_logic_vector(to_unsigned( 245,8)),
			14521 => std_logic_vector(to_unsigned( 226,8)),
			14522 => std_logic_vector(to_unsigned( 87,8)),
			14523 => std_logic_vector(to_unsigned( 26,8)),
			14524 => std_logic_vector(to_unsigned( 107,8)),
			14525 => std_logic_vector(to_unsigned( 150,8)),
			14526 => std_logic_vector(to_unsigned( 140,8)),
			14527 => std_logic_vector(to_unsigned( 124,8)),
			14528 => std_logic_vector(to_unsigned( 213,8)),
			14529 => std_logic_vector(to_unsigned( 164,8)),
			14530 => std_logic_vector(to_unsigned( 140,8)),
			14531 => std_logic_vector(to_unsigned( 34,8)),
			14532 => std_logic_vector(to_unsigned( 1,8)),
			14533 => std_logic_vector(to_unsigned( 174,8)),
			14534 => std_logic_vector(to_unsigned( 204,8)),
			14535 => std_logic_vector(to_unsigned( 229,8)),
			14536 => std_logic_vector(to_unsigned( 107,8)),
			14537 => std_logic_vector(to_unsigned( 100,8)),
			14538 => std_logic_vector(to_unsigned( 82,8)),
			14539 => std_logic_vector(to_unsigned( 251,8)),
			14540 => std_logic_vector(to_unsigned( 230,8)),
			14541 => std_logic_vector(to_unsigned( 190,8)),
			14542 => std_logic_vector(to_unsigned( 128,8)),
			14543 => std_logic_vector(to_unsigned( 145,8)),
			14544 => std_logic_vector(to_unsigned( 196,8)),
			14545 => std_logic_vector(to_unsigned( 134,8)),
			14546 => std_logic_vector(to_unsigned( 84,8)),
			14547 => std_logic_vector(to_unsigned( 235,8)),
			14548 => std_logic_vector(to_unsigned( 17,8)),
			14549 => std_logic_vector(to_unsigned( 129,8)),
			14550 => std_logic_vector(to_unsigned( 195,8)),
			14551 => std_logic_vector(to_unsigned( 180,8)),
			14552 => std_logic_vector(to_unsigned( 120,8)),
			14553 => std_logic_vector(to_unsigned( 7,8)),
			14554 => std_logic_vector(to_unsigned( 38,8)),
			14555 => std_logic_vector(to_unsigned( 62,8)),
			14556 => std_logic_vector(to_unsigned( 213,8)),
			14557 => std_logic_vector(to_unsigned( 88,8)),
			14558 => std_logic_vector(to_unsigned( 89,8)),
			14559 => std_logic_vector(to_unsigned( 253,8)),
			14560 => std_logic_vector(to_unsigned( 169,8)),
			14561 => std_logic_vector(to_unsigned( 231,8)),
			14562 => std_logic_vector(to_unsigned( 75,8)),
			14563 => std_logic_vector(to_unsigned( 191,8)),
			14564 => std_logic_vector(to_unsigned( 172,8)),
			14565 => std_logic_vector(to_unsigned( 119,8)),
			14566 => std_logic_vector(to_unsigned( 206,8)),
			14567 => std_logic_vector(to_unsigned( 157,8)),
			14568 => std_logic_vector(to_unsigned( 6,8)),
			14569 => std_logic_vector(to_unsigned( 210,8)),
			14570 => std_logic_vector(to_unsigned( 110,8)),
			14571 => std_logic_vector(to_unsigned( 223,8)),
			14572 => std_logic_vector(to_unsigned( 128,8)),
			14573 => std_logic_vector(to_unsigned( 47,8)),
			14574 => std_logic_vector(to_unsigned( 156,8)),
			14575 => std_logic_vector(to_unsigned( 100,8)),
			14576 => std_logic_vector(to_unsigned( 243,8)),
			14577 => std_logic_vector(to_unsigned( 140,8)),
			14578 => std_logic_vector(to_unsigned( 94,8)),
			14579 => std_logic_vector(to_unsigned( 68,8)),
			14580 => std_logic_vector(to_unsigned( 247,8)),
			14581 => std_logic_vector(to_unsigned( 243,8)),
			14582 => std_logic_vector(to_unsigned( 26,8)),
			14583 => std_logic_vector(to_unsigned( 213,8)),
			14584 => std_logic_vector(to_unsigned( 253,8)),
			14585 => std_logic_vector(to_unsigned( 21,8)),
			14586 => std_logic_vector(to_unsigned( 78,8)),
			14587 => std_logic_vector(to_unsigned( 1,8)),
			14588 => std_logic_vector(to_unsigned( 48,8)),
			14589 => std_logic_vector(to_unsigned( 27,8)),
			14590 => std_logic_vector(to_unsigned( 20,8)),
			14591 => std_logic_vector(to_unsigned( 224,8)),
			14592 => std_logic_vector(to_unsigned( 212,8)),
			14593 => std_logic_vector(to_unsigned( 11,8)),
			14594 => std_logic_vector(to_unsigned( 168,8)),
			14595 => std_logic_vector(to_unsigned( 6,8)),
			14596 => std_logic_vector(to_unsigned( 109,8)),
			14597 => std_logic_vector(to_unsigned( 174,8)),
			14598 => std_logic_vector(to_unsigned( 91,8)),
			14599 => std_logic_vector(to_unsigned( 62,8)),
			14600 => std_logic_vector(to_unsigned( 234,8)),
			14601 => std_logic_vector(to_unsigned( 53,8)),
			14602 => std_logic_vector(to_unsigned( 20,8)),
			14603 => std_logic_vector(to_unsigned( 75,8)),
			14604 => std_logic_vector(to_unsigned( 153,8)),
			14605 => std_logic_vector(to_unsigned( 186,8)),
			14606 => std_logic_vector(to_unsigned( 24,8)),
			14607 => std_logic_vector(to_unsigned( 221,8)),
			14608 => std_logic_vector(to_unsigned( 188,8)),
			14609 => std_logic_vector(to_unsigned( 233,8)),
			14610 => std_logic_vector(to_unsigned( 27,8)),
			14611 => std_logic_vector(to_unsigned( 150,8)),
			14612 => std_logic_vector(to_unsigned( 28,8)),
			14613 => std_logic_vector(to_unsigned( 7,8)),
			14614 => std_logic_vector(to_unsigned( 22,8)),
			14615 => std_logic_vector(to_unsigned( 161,8)),
			14616 => std_logic_vector(to_unsigned( 204,8)),
			14617 => std_logic_vector(to_unsigned( 121,8)),
			14618 => std_logic_vector(to_unsigned( 209,8)),
			14619 => std_logic_vector(to_unsigned( 184,8)),
			14620 => std_logic_vector(to_unsigned( 137,8)),
			14621 => std_logic_vector(to_unsigned( 76,8)),
			14622 => std_logic_vector(to_unsigned( 211,8)),
			14623 => std_logic_vector(to_unsigned( 200,8)),
			14624 => std_logic_vector(to_unsigned( 137,8)),
			14625 => std_logic_vector(to_unsigned( 71,8)),
			14626 => std_logic_vector(to_unsigned( 247,8)),
			14627 => std_logic_vector(to_unsigned( 212,8)),
			14628 => std_logic_vector(to_unsigned( 200,8)),
			14629 => std_logic_vector(to_unsigned( 111,8)),
			14630 => std_logic_vector(to_unsigned( 203,8)),
			14631 => std_logic_vector(to_unsigned( 40,8)),
			14632 => std_logic_vector(to_unsigned( 207,8)),
			14633 => std_logic_vector(to_unsigned( 255,8)),
			14634 => std_logic_vector(to_unsigned( 132,8)),
			14635 => std_logic_vector(to_unsigned( 232,8)),
			14636 => std_logic_vector(to_unsigned( 81,8)),
			14637 => std_logic_vector(to_unsigned( 100,8)),
			14638 => std_logic_vector(to_unsigned( 174,8)),
			14639 => std_logic_vector(to_unsigned( 27,8)),
			14640 => std_logic_vector(to_unsigned( 145,8)),
			14641 => std_logic_vector(to_unsigned( 199,8)),
			14642 => std_logic_vector(to_unsigned( 99,8)),
			14643 => std_logic_vector(to_unsigned( 237,8)),
			14644 => std_logic_vector(to_unsigned( 129,8)),
			14645 => std_logic_vector(to_unsigned( 83,8)),
			14646 => std_logic_vector(to_unsigned( 1,8)),
			14647 => std_logic_vector(to_unsigned( 129,8)),
			14648 => std_logic_vector(to_unsigned( 40,8)),
			14649 => std_logic_vector(to_unsigned( 220,8)),
			14650 => std_logic_vector(to_unsigned( 126,8)),
			14651 => std_logic_vector(to_unsigned( 95,8)),
			14652 => std_logic_vector(to_unsigned( 233,8)),
			14653 => std_logic_vector(to_unsigned( 215,8)),
			14654 => std_logic_vector(to_unsigned( 131,8)),
			14655 => std_logic_vector(to_unsigned( 61,8)),
			14656 => std_logic_vector(to_unsigned( 133,8)),
			14657 => std_logic_vector(to_unsigned( 232,8)),
			14658 => std_logic_vector(to_unsigned( 86,8)),
			14659 => std_logic_vector(to_unsigned( 16,8)),
			14660 => std_logic_vector(to_unsigned( 118,8)),
			14661 => std_logic_vector(to_unsigned( 199,8)),
			14662 => std_logic_vector(to_unsigned( 238,8)),
			14663 => std_logic_vector(to_unsigned( 152,8)),
			14664 => std_logic_vector(to_unsigned( 76,8)),
			14665 => std_logic_vector(to_unsigned( 176,8)),
			14666 => std_logic_vector(to_unsigned( 203,8)),
			14667 => std_logic_vector(to_unsigned( 159,8)),
			14668 => std_logic_vector(to_unsigned( 199,8)),
			14669 => std_logic_vector(to_unsigned( 210,8)),
			14670 => std_logic_vector(to_unsigned( 210,8)),
			14671 => std_logic_vector(to_unsigned( 175,8)),
			14672 => std_logic_vector(to_unsigned( 145,8)),
			14673 => std_logic_vector(to_unsigned( 116,8)),
			14674 => std_logic_vector(to_unsigned( 49,8)),
			14675 => std_logic_vector(to_unsigned( 212,8)),
			14676 => std_logic_vector(to_unsigned( 157,8)),
			14677 => std_logic_vector(to_unsigned( 5,8)),
			14678 => std_logic_vector(to_unsigned( 208,8)),
			14679 => std_logic_vector(to_unsigned( 81,8)),
			14680 => std_logic_vector(to_unsigned( 249,8)),
			14681 => std_logic_vector(to_unsigned( 140,8)),
			14682 => std_logic_vector(to_unsigned( 86,8)),
			14683 => std_logic_vector(to_unsigned( 126,8)),
			14684 => std_logic_vector(to_unsigned( 62,8)),
			14685 => std_logic_vector(to_unsigned( 193,8)),
			14686 => std_logic_vector(to_unsigned( 241,8)),
			14687 => std_logic_vector(to_unsigned( 88,8)),
			14688 => std_logic_vector(to_unsigned( 6,8)),
			14689 => std_logic_vector(to_unsigned( 180,8)),
			14690 => std_logic_vector(to_unsigned( 52,8)),
			14691 => std_logic_vector(to_unsigned( 214,8)),
			14692 => std_logic_vector(to_unsigned( 195,8)),
			14693 => std_logic_vector(to_unsigned( 231,8)),
			14694 => std_logic_vector(to_unsigned( 15,8)),
			14695 => std_logic_vector(to_unsigned( 226,8)),
			14696 => std_logic_vector(to_unsigned( 12,8)),
			14697 => std_logic_vector(to_unsigned( 192,8)),
			14698 => std_logic_vector(to_unsigned( 93,8)),
			14699 => std_logic_vector(to_unsigned( 164,8)),
			14700 => std_logic_vector(to_unsigned( 250,8)),
			14701 => std_logic_vector(to_unsigned( 63,8)),
			14702 => std_logic_vector(to_unsigned( 197,8)),
			14703 => std_logic_vector(to_unsigned( 131,8)),
			14704 => std_logic_vector(to_unsigned( 117,8)),
			14705 => std_logic_vector(to_unsigned( 75,8)),
			14706 => std_logic_vector(to_unsigned( 191,8)),
			14707 => std_logic_vector(to_unsigned( 224,8)),
			14708 => std_logic_vector(to_unsigned( 234,8)),
			14709 => std_logic_vector(to_unsigned( 209,8)),
			14710 => std_logic_vector(to_unsigned( 20,8)),
			14711 => std_logic_vector(to_unsigned( 34,8)),
			14712 => std_logic_vector(to_unsigned( 77,8)),
			14713 => std_logic_vector(to_unsigned( 209,8)),
			14714 => std_logic_vector(to_unsigned( 77,8)),
			14715 => std_logic_vector(to_unsigned( 30,8)),
			14716 => std_logic_vector(to_unsigned( 162,8)),
			14717 => std_logic_vector(to_unsigned( 145,8)),
			14718 => std_logic_vector(to_unsigned( 149,8)),
			14719 => std_logic_vector(to_unsigned( 224,8)),
			14720 => std_logic_vector(to_unsigned( 27,8)),
			14721 => std_logic_vector(to_unsigned( 155,8)),
			14722 => std_logic_vector(to_unsigned( 54,8)),
			14723 => std_logic_vector(to_unsigned( 80,8)),
			14724 => std_logic_vector(to_unsigned( 186,8)),
			14725 => std_logic_vector(to_unsigned( 16,8)),
			14726 => std_logic_vector(to_unsigned( 77,8)),
			14727 => std_logic_vector(to_unsigned( 51,8)),
			14728 => std_logic_vector(to_unsigned( 146,8)),
			14729 => std_logic_vector(to_unsigned( 53,8)),
			14730 => std_logic_vector(to_unsigned( 127,8)),
			14731 => std_logic_vector(to_unsigned( 152,8)),
			14732 => std_logic_vector(to_unsigned( 131,8)),
			14733 => std_logic_vector(to_unsigned( 60,8)),
			14734 => std_logic_vector(to_unsigned( 165,8)),
			14735 => std_logic_vector(to_unsigned( 178,8)),
			14736 => std_logic_vector(to_unsigned( 11,8)),
			14737 => std_logic_vector(to_unsigned( 55,8)),
			14738 => std_logic_vector(to_unsigned( 121,8)),
			14739 => std_logic_vector(to_unsigned( 71,8)),
			14740 => std_logic_vector(to_unsigned( 119,8)),
			14741 => std_logic_vector(to_unsigned( 194,8)),
			14742 => std_logic_vector(to_unsigned( 141,8)),
			14743 => std_logic_vector(to_unsigned( 230,8)),
			14744 => std_logic_vector(to_unsigned( 223,8)),
			14745 => std_logic_vector(to_unsigned( 201,8)),
			14746 => std_logic_vector(to_unsigned( 211,8)),
			14747 => std_logic_vector(to_unsigned( 171,8)),
			14748 => std_logic_vector(to_unsigned( 234,8)),
			14749 => std_logic_vector(to_unsigned( 143,8)),
			14750 => std_logic_vector(to_unsigned( 98,8)),
			14751 => std_logic_vector(to_unsigned( 255,8)),
			14752 => std_logic_vector(to_unsigned( 130,8)),
			14753 => std_logic_vector(to_unsigned( 137,8)),
			14754 => std_logic_vector(to_unsigned( 104,8)),
			14755 => std_logic_vector(to_unsigned( 200,8)),
			14756 => std_logic_vector(to_unsigned( 15,8)),
			14757 => std_logic_vector(to_unsigned( 170,8)),
			14758 => std_logic_vector(to_unsigned( 30,8)),
			14759 => std_logic_vector(to_unsigned( 255,8)),
			14760 => std_logic_vector(to_unsigned( 251,8)),
			14761 => std_logic_vector(to_unsigned( 210,8)),
			14762 => std_logic_vector(to_unsigned( 248,8)),
			14763 => std_logic_vector(to_unsigned( 75,8)),
			14764 => std_logic_vector(to_unsigned( 87,8)),
			14765 => std_logic_vector(to_unsigned( 212,8)),
			14766 => std_logic_vector(to_unsigned( 88,8)),
			14767 => std_logic_vector(to_unsigned( 188,8)),
			14768 => std_logic_vector(to_unsigned( 167,8)),
			14769 => std_logic_vector(to_unsigned( 31,8)),
			14770 => std_logic_vector(to_unsigned( 89,8)),
			14771 => std_logic_vector(to_unsigned( 204,8)),
			14772 => std_logic_vector(to_unsigned( 24,8)),
			14773 => std_logic_vector(to_unsigned( 90,8)),
			14774 => std_logic_vector(to_unsigned( 71,8)),
			14775 => std_logic_vector(to_unsigned( 23,8)),
			14776 => std_logic_vector(to_unsigned( 248,8)),
			14777 => std_logic_vector(to_unsigned( 80,8)),
			14778 => std_logic_vector(to_unsigned( 90,8)),
			14779 => std_logic_vector(to_unsigned( 123,8)),
			14780 => std_logic_vector(to_unsigned( 179,8)),
			14781 => std_logic_vector(to_unsigned( 176,8)),
			14782 => std_logic_vector(to_unsigned( 85,8)),
			14783 => std_logic_vector(to_unsigned( 236,8)),
			14784 => std_logic_vector(to_unsigned( 41,8)),
			14785 => std_logic_vector(to_unsigned( 34,8)),
			14786 => std_logic_vector(to_unsigned( 152,8)),
			14787 => std_logic_vector(to_unsigned( 58,8)),
			14788 => std_logic_vector(to_unsigned( 136,8)),
			14789 => std_logic_vector(to_unsigned( 34,8)),
			14790 => std_logic_vector(to_unsigned( 96,8)),
			14791 => std_logic_vector(to_unsigned( 150,8)),
			14792 => std_logic_vector(to_unsigned( 250,8)),
			14793 => std_logic_vector(to_unsigned( 224,8)),
			14794 => std_logic_vector(to_unsigned( 166,8)),
			14795 => std_logic_vector(to_unsigned( 166,8)),
			14796 => std_logic_vector(to_unsigned( 214,8)),
			14797 => std_logic_vector(to_unsigned( 148,8)),
			14798 => std_logic_vector(to_unsigned( 144,8)),
			14799 => std_logic_vector(to_unsigned( 127,8)),
			14800 => std_logic_vector(to_unsigned( 112,8)),
			14801 => std_logic_vector(to_unsigned( 116,8)),
			14802 => std_logic_vector(to_unsigned( 132,8)),
			14803 => std_logic_vector(to_unsigned( 244,8)),
			14804 => std_logic_vector(to_unsigned( 69,8)),
			14805 => std_logic_vector(to_unsigned( 174,8)),
			14806 => std_logic_vector(to_unsigned( 11,8)),
			14807 => std_logic_vector(to_unsigned( 209,8)),
			14808 => std_logic_vector(to_unsigned( 241,8)),
			14809 => std_logic_vector(to_unsigned( 214,8)),
			14810 => std_logic_vector(to_unsigned( 223,8)),
			14811 => std_logic_vector(to_unsigned( 9,8)),
			14812 => std_logic_vector(to_unsigned( 131,8)),
			14813 => std_logic_vector(to_unsigned( 56,8)),
			14814 => std_logic_vector(to_unsigned( 204,8)),
			14815 => std_logic_vector(to_unsigned( 102,8)),
			14816 => std_logic_vector(to_unsigned( 7,8)),
			14817 => std_logic_vector(to_unsigned( 87,8)),
			14818 => std_logic_vector(to_unsigned( 96,8)),
			14819 => std_logic_vector(to_unsigned( 213,8)),
			14820 => std_logic_vector(to_unsigned( 220,8)),
			14821 => std_logic_vector(to_unsigned( 102,8)),
			14822 => std_logic_vector(to_unsigned( 146,8)),
			14823 => std_logic_vector(to_unsigned( 97,8)),
			14824 => std_logic_vector(to_unsigned( 246,8)),
			14825 => std_logic_vector(to_unsigned( 254,8)),
			14826 => std_logic_vector(to_unsigned( 36,8)),
			14827 => std_logic_vector(to_unsigned( 29,8)),
			14828 => std_logic_vector(to_unsigned( 68,8)),
			14829 => std_logic_vector(to_unsigned( 178,8)),
			14830 => std_logic_vector(to_unsigned( 106,8)),
			14831 => std_logic_vector(to_unsigned( 16,8)),
			14832 => std_logic_vector(to_unsigned( 237,8)),
			14833 => std_logic_vector(to_unsigned( 7,8)),
			14834 => std_logic_vector(to_unsigned( 99,8)),
			14835 => std_logic_vector(to_unsigned( 181,8)),
			14836 => std_logic_vector(to_unsigned( 145,8)),
			14837 => std_logic_vector(to_unsigned( 188,8)),
			14838 => std_logic_vector(to_unsigned( 207,8)),
			14839 => std_logic_vector(to_unsigned( 98,8)),
			14840 => std_logic_vector(to_unsigned( 220,8)),
			14841 => std_logic_vector(to_unsigned( 233,8)),
			14842 => std_logic_vector(to_unsigned( 103,8)),
			14843 => std_logic_vector(to_unsigned( 247,8)),
			14844 => std_logic_vector(to_unsigned( 17,8)),
			14845 => std_logic_vector(to_unsigned( 68,8)),
			14846 => std_logic_vector(to_unsigned( 13,8)),
			14847 => std_logic_vector(to_unsigned( 143,8)),
			14848 => std_logic_vector(to_unsigned( 201,8)),
			14849 => std_logic_vector(to_unsigned( 136,8)),
			14850 => std_logic_vector(to_unsigned( 154,8)),
			14851 => std_logic_vector(to_unsigned( 145,8)),
			14852 => std_logic_vector(to_unsigned( 159,8)),
			14853 => std_logic_vector(to_unsigned( 223,8)),
			14854 => std_logic_vector(to_unsigned( 100,8)),
			14855 => std_logic_vector(to_unsigned( 132,8)),
			14856 => std_logic_vector(to_unsigned( 227,8)),
			14857 => std_logic_vector(to_unsigned( 73,8)),
			14858 => std_logic_vector(to_unsigned( 52,8)),
			14859 => std_logic_vector(to_unsigned( 141,8)),
			14860 => std_logic_vector(to_unsigned( 70,8)),
			14861 => std_logic_vector(to_unsigned( 6,8)),
			14862 => std_logic_vector(to_unsigned( 125,8)),
			14863 => std_logic_vector(to_unsigned( 143,8)),
			14864 => std_logic_vector(to_unsigned( 64,8)),
			14865 => std_logic_vector(to_unsigned( 219,8)),
			14866 => std_logic_vector(to_unsigned( 170,8)),
			14867 => std_logic_vector(to_unsigned( 11,8)),
			14868 => std_logic_vector(to_unsigned( 180,8)),
			14869 => std_logic_vector(to_unsigned( 26,8)),
			14870 => std_logic_vector(to_unsigned( 13,8)),
			14871 => std_logic_vector(to_unsigned( 166,8)),
			14872 => std_logic_vector(to_unsigned( 76,8)),
			14873 => std_logic_vector(to_unsigned( 227,8)),
			14874 => std_logic_vector(to_unsigned( 122,8)),
			14875 => std_logic_vector(to_unsigned( 5,8)),
			14876 => std_logic_vector(to_unsigned( 143,8)),
			14877 => std_logic_vector(to_unsigned( 154,8)),
			14878 => std_logic_vector(to_unsigned( 24,8)),
			14879 => std_logic_vector(to_unsigned( 163,8)),
			14880 => std_logic_vector(to_unsigned( 23,8)),
			14881 => std_logic_vector(to_unsigned( 165,8)),
			14882 => std_logic_vector(to_unsigned( 140,8)),
			14883 => std_logic_vector(to_unsigned( 37,8)),
			14884 => std_logic_vector(to_unsigned( 24,8)),
			14885 => std_logic_vector(to_unsigned( 55,8)),
			14886 => std_logic_vector(to_unsigned( 43,8)),
			14887 => std_logic_vector(to_unsigned( 95,8)),
			14888 => std_logic_vector(to_unsigned( 149,8)),
			14889 => std_logic_vector(to_unsigned( 226,8)),
			14890 => std_logic_vector(to_unsigned( 161,8)),
			14891 => std_logic_vector(to_unsigned( 122,8)),
			14892 => std_logic_vector(to_unsigned( 99,8)),
			14893 => std_logic_vector(to_unsigned( 201,8)),
			14894 => std_logic_vector(to_unsigned( 14,8)),
			14895 => std_logic_vector(to_unsigned( 182,8)),
			14896 => std_logic_vector(to_unsigned( 135,8)),
			14897 => std_logic_vector(to_unsigned( 179,8)),
			14898 => std_logic_vector(to_unsigned( 10,8)),
			14899 => std_logic_vector(to_unsigned( 53,8)),
			14900 => std_logic_vector(to_unsigned( 22,8)),
			14901 => std_logic_vector(to_unsigned( 226,8)),
			14902 => std_logic_vector(to_unsigned( 82,8)),
			14903 => std_logic_vector(to_unsigned( 226,8)),
			14904 => std_logic_vector(to_unsigned( 8,8)),
			14905 => std_logic_vector(to_unsigned( 63,8)),
			14906 => std_logic_vector(to_unsigned( 182,8)),
			14907 => std_logic_vector(to_unsigned( 95,8)),
			14908 => std_logic_vector(to_unsigned( 129,8)),
			14909 => std_logic_vector(to_unsigned( 111,8)),
			14910 => std_logic_vector(to_unsigned( 68,8)),
			14911 => std_logic_vector(to_unsigned( 217,8)),
			14912 => std_logic_vector(to_unsigned( 113,8)),
			14913 => std_logic_vector(to_unsigned( 20,8)),
			14914 => std_logic_vector(to_unsigned( 48,8)),
			14915 => std_logic_vector(to_unsigned( 90,8)),
			14916 => std_logic_vector(to_unsigned( 44,8)),
			14917 => std_logic_vector(to_unsigned( 38,8)),
			14918 => std_logic_vector(to_unsigned( 58,8)),
			14919 => std_logic_vector(to_unsigned( 213,8)),
			14920 => std_logic_vector(to_unsigned( 26,8)),
			14921 => std_logic_vector(to_unsigned( 232,8)),
			14922 => std_logic_vector(to_unsigned( 40,8)),
			14923 => std_logic_vector(to_unsigned( 222,8)),
			14924 => std_logic_vector(to_unsigned( 118,8)),
			14925 => std_logic_vector(to_unsigned( 150,8)),
			14926 => std_logic_vector(to_unsigned( 63,8)),
			14927 => std_logic_vector(to_unsigned( 159,8)),
			14928 => std_logic_vector(to_unsigned( 158,8)),
			14929 => std_logic_vector(to_unsigned( 54,8)),
			14930 => std_logic_vector(to_unsigned( 254,8)),
			14931 => std_logic_vector(to_unsigned( 151,8)),
			14932 => std_logic_vector(to_unsigned( 51,8)),
			14933 => std_logic_vector(to_unsigned( 238,8)),
			14934 => std_logic_vector(to_unsigned( 184,8)),
			14935 => std_logic_vector(to_unsigned( 32,8)),
			14936 => std_logic_vector(to_unsigned( 99,8)),
			14937 => std_logic_vector(to_unsigned( 242,8)),
			14938 => std_logic_vector(to_unsigned( 228,8)),
			14939 => std_logic_vector(to_unsigned( 241,8)),
			14940 => std_logic_vector(to_unsigned( 252,8)),
			14941 => std_logic_vector(to_unsigned( 156,8)),
			14942 => std_logic_vector(to_unsigned( 243,8)),
			14943 => std_logic_vector(to_unsigned( 246,8)),
			14944 => std_logic_vector(to_unsigned( 216,8)),
			14945 => std_logic_vector(to_unsigned( 86,8)),
			14946 => std_logic_vector(to_unsigned( 239,8)),
			14947 => std_logic_vector(to_unsigned( 83,8)),
			14948 => std_logic_vector(to_unsigned( 36,8)),
			14949 => std_logic_vector(to_unsigned( 95,8)),
			14950 => std_logic_vector(to_unsigned( 5,8)),
			14951 => std_logic_vector(to_unsigned( 76,8)),
			14952 => std_logic_vector(to_unsigned( 199,8)),
			14953 => std_logic_vector(to_unsigned( 50,8)),
			14954 => std_logic_vector(to_unsigned( 15,8)),
			14955 => std_logic_vector(to_unsigned( 44,8)),
			14956 => std_logic_vector(to_unsigned( 113,8)),
			14957 => std_logic_vector(to_unsigned( 190,8)),
			14958 => std_logic_vector(to_unsigned( 43,8)),
			14959 => std_logic_vector(to_unsigned( 210,8)),
			14960 => std_logic_vector(to_unsigned( 67,8)),
			14961 => std_logic_vector(to_unsigned( 187,8)),
			14962 => std_logic_vector(to_unsigned( 168,8)),
			14963 => std_logic_vector(to_unsigned( 11,8)),
			14964 => std_logic_vector(to_unsigned( 96,8)),
			14965 => std_logic_vector(to_unsigned( 209,8)),
			14966 => std_logic_vector(to_unsigned( 213,8)),
			14967 => std_logic_vector(to_unsigned( 165,8)),
			14968 => std_logic_vector(to_unsigned( 124,8)),
			14969 => std_logic_vector(to_unsigned( 124,8)),
			14970 => std_logic_vector(to_unsigned( 35,8)),
			14971 => std_logic_vector(to_unsigned( 96,8)),
			14972 => std_logic_vector(to_unsigned( 100,8)),
			14973 => std_logic_vector(to_unsigned( 103,8)),
			14974 => std_logic_vector(to_unsigned( 65,8)),
			14975 => std_logic_vector(to_unsigned( 119,8)),
			14976 => std_logic_vector(to_unsigned( 226,8)),
			14977 => std_logic_vector(to_unsigned( 229,8)),
			14978 => std_logic_vector(to_unsigned( 200,8)),
			14979 => std_logic_vector(to_unsigned( 134,8)),
			14980 => std_logic_vector(to_unsigned( 110,8)),
			14981 => std_logic_vector(to_unsigned( 231,8)),
			14982 => std_logic_vector(to_unsigned( 158,8)),
			14983 => std_logic_vector(to_unsigned( 137,8)),
			14984 => std_logic_vector(to_unsigned( 185,8)),
			14985 => std_logic_vector(to_unsigned( 210,8)),
			14986 => std_logic_vector(to_unsigned( 72,8)),
			14987 => std_logic_vector(to_unsigned( 199,8)),
			14988 => std_logic_vector(to_unsigned( 234,8)),
			14989 => std_logic_vector(to_unsigned( 204,8)),
			14990 => std_logic_vector(to_unsigned( 122,8)),
			14991 => std_logic_vector(to_unsigned( 160,8)),
			14992 => std_logic_vector(to_unsigned( 114,8)),
			14993 => std_logic_vector(to_unsigned( 89,8)),
			14994 => std_logic_vector(to_unsigned( 160,8)),
			14995 => std_logic_vector(to_unsigned( 104,8)),
			14996 => std_logic_vector(to_unsigned( 125,8)),
			14997 => std_logic_vector(to_unsigned( 242,8)),
			14998 => std_logic_vector(to_unsigned( 3,8)),
			14999 => std_logic_vector(to_unsigned( 150,8)),
			15000 => std_logic_vector(to_unsigned( 139,8)),
			15001 => std_logic_vector(to_unsigned( 225,8)),
			15002 => std_logic_vector(to_unsigned( 12,8)),
			15003 => std_logic_vector(to_unsigned( 220,8)),
			15004 => std_logic_vector(to_unsigned( 107,8)),
			15005 => std_logic_vector(to_unsigned( 142,8)),
			15006 => std_logic_vector(to_unsigned( 31,8)),
			15007 => std_logic_vector(to_unsigned( 192,8)),
			15008 => std_logic_vector(to_unsigned( 177,8)),
			15009 => std_logic_vector(to_unsigned( 49,8)),
			15010 => std_logic_vector(to_unsigned( 9,8)),
			15011 => std_logic_vector(to_unsigned( 192,8)),
			15012 => std_logic_vector(to_unsigned( 155,8)),
			15013 => std_logic_vector(to_unsigned( 91,8)),
			15014 => std_logic_vector(to_unsigned( 173,8)),
			15015 => std_logic_vector(to_unsigned( 29,8)),
			15016 => std_logic_vector(to_unsigned( 127,8)),
			15017 => std_logic_vector(to_unsigned( 125,8)),
			15018 => std_logic_vector(to_unsigned( 102,8)),
			15019 => std_logic_vector(to_unsigned( 115,8)),
			15020 => std_logic_vector(to_unsigned( 123,8)),
			15021 => std_logic_vector(to_unsigned( 228,8)),
			15022 => std_logic_vector(to_unsigned( 3,8)),
			15023 => std_logic_vector(to_unsigned( 48,8)),
			15024 => std_logic_vector(to_unsigned( 247,8)),
			15025 => std_logic_vector(to_unsigned( 130,8)),
			15026 => std_logic_vector(to_unsigned( 253,8)),
			15027 => std_logic_vector(to_unsigned( 113,8)),
			15028 => std_logic_vector(to_unsigned( 166,8)),
			15029 => std_logic_vector(to_unsigned( 41,8)),
			15030 => std_logic_vector(to_unsigned( 251,8)),
			15031 => std_logic_vector(to_unsigned( 52,8)),
			15032 => std_logic_vector(to_unsigned( 186,8)),
			15033 => std_logic_vector(to_unsigned( 84,8)),
			15034 => std_logic_vector(to_unsigned( 23,8)),
			15035 => std_logic_vector(to_unsigned( 223,8)),
			15036 => std_logic_vector(to_unsigned( 15,8)),
			15037 => std_logic_vector(to_unsigned( 105,8)),
			15038 => std_logic_vector(to_unsigned( 52,8)),
			15039 => std_logic_vector(to_unsigned( 39,8)),
			15040 => std_logic_vector(to_unsigned( 142,8)),
			15041 => std_logic_vector(to_unsigned( 6,8)),
			15042 => std_logic_vector(to_unsigned( 196,8)),
			15043 => std_logic_vector(to_unsigned( 146,8)),
			15044 => std_logic_vector(to_unsigned( 86,8)),
			15045 => std_logic_vector(to_unsigned( 138,8)),
			15046 => std_logic_vector(to_unsigned( 230,8)),
			15047 => std_logic_vector(to_unsigned( 249,8)),
			15048 => std_logic_vector(to_unsigned( 107,8)),
			15049 => std_logic_vector(to_unsigned( 143,8)),
			15050 => std_logic_vector(to_unsigned( 232,8)),
			15051 => std_logic_vector(to_unsigned( 126,8)),
			15052 => std_logic_vector(to_unsigned( 109,8)),
			15053 => std_logic_vector(to_unsigned( 211,8)),
			15054 => std_logic_vector(to_unsigned( 255,8)),
			15055 => std_logic_vector(to_unsigned( 194,8)),
			15056 => std_logic_vector(to_unsigned( 226,8)),
			15057 => std_logic_vector(to_unsigned( 88,8)),
			15058 => std_logic_vector(to_unsigned( 185,8)),
			15059 => std_logic_vector(to_unsigned( 202,8)),
			15060 => std_logic_vector(to_unsigned( 182,8)),
			15061 => std_logic_vector(to_unsigned( 147,8)),
			15062 => std_logic_vector(to_unsigned( 115,8)),
			15063 => std_logic_vector(to_unsigned( 109,8)),
			15064 => std_logic_vector(to_unsigned( 225,8)),
			15065 => std_logic_vector(to_unsigned( 97,8)),
			15066 => std_logic_vector(to_unsigned( 65,8)),
			15067 => std_logic_vector(to_unsigned( 121,8)),
			15068 => std_logic_vector(to_unsigned( 181,8)),
			15069 => std_logic_vector(to_unsigned( 61,8)),
			15070 => std_logic_vector(to_unsigned( 135,8)),
			15071 => std_logic_vector(to_unsigned( 88,8)),
			15072 => std_logic_vector(to_unsigned( 85,8)),
			15073 => std_logic_vector(to_unsigned( 188,8)),
			15074 => std_logic_vector(to_unsigned( 109,8)),
			15075 => std_logic_vector(to_unsigned( 181,8)),
			15076 => std_logic_vector(to_unsigned( 187,8)),
			15077 => std_logic_vector(to_unsigned( 249,8)),
			15078 => std_logic_vector(to_unsigned( 124,8)),
			15079 => std_logic_vector(to_unsigned( 159,8)),
			15080 => std_logic_vector(to_unsigned( 15,8)),
			15081 => std_logic_vector(to_unsigned( 159,8)),
			15082 => std_logic_vector(to_unsigned( 115,8)),
			15083 => std_logic_vector(to_unsigned( 154,8)),
			15084 => std_logic_vector(to_unsigned( 168,8)),
			15085 => std_logic_vector(to_unsigned( 90,8)),
			15086 => std_logic_vector(to_unsigned( 180,8)),
			15087 => std_logic_vector(to_unsigned( 231,8)),
			15088 => std_logic_vector(to_unsigned( 168,8)),
			15089 => std_logic_vector(to_unsigned( 245,8)),
			15090 => std_logic_vector(to_unsigned( 117,8)),
			15091 => std_logic_vector(to_unsigned( 165,8)),
			15092 => std_logic_vector(to_unsigned( 88,8)),
			15093 => std_logic_vector(to_unsigned( 148,8)),
			15094 => std_logic_vector(to_unsigned( 216,8)),
			15095 => std_logic_vector(to_unsigned( 75,8)),
			15096 => std_logic_vector(to_unsigned( 228,8)),
			15097 => std_logic_vector(to_unsigned( 55,8)),
			15098 => std_logic_vector(to_unsigned( 169,8)),
			15099 => std_logic_vector(to_unsigned( 64,8)),
			15100 => std_logic_vector(to_unsigned( 23,8)),
			15101 => std_logic_vector(to_unsigned( 97,8)),
			15102 => std_logic_vector(to_unsigned( 69,8)),
			15103 => std_logic_vector(to_unsigned( 167,8)),
			15104 => std_logic_vector(to_unsigned( 169,8)),
			15105 => std_logic_vector(to_unsigned( 69,8)),
			15106 => std_logic_vector(to_unsigned( 162,8)),
			15107 => std_logic_vector(to_unsigned( 163,8)),
			15108 => std_logic_vector(to_unsigned( 172,8)),
			15109 => std_logic_vector(to_unsigned( 129,8)),
			15110 => std_logic_vector(to_unsigned( 201,8)),
			15111 => std_logic_vector(to_unsigned( 77,8)),
			15112 => std_logic_vector(to_unsigned( 71,8)),
			15113 => std_logic_vector(to_unsigned( 22,8)),
			15114 => std_logic_vector(to_unsigned( 237,8)),
			15115 => std_logic_vector(to_unsigned( 46,8)),
			15116 => std_logic_vector(to_unsigned( 85,8)),
			15117 => std_logic_vector(to_unsigned( 217,8)),
			15118 => std_logic_vector(to_unsigned( 17,8)),
			15119 => std_logic_vector(to_unsigned( 185,8)),
			15120 => std_logic_vector(to_unsigned( 80,8)),
			15121 => std_logic_vector(to_unsigned( 79,8)),
			15122 => std_logic_vector(to_unsigned( 104,8)),
			15123 => std_logic_vector(to_unsigned( 20,8)),
			15124 => std_logic_vector(to_unsigned( 107,8)),
			15125 => std_logic_vector(to_unsigned( 156,8)),
			15126 => std_logic_vector(to_unsigned( 112,8)),
			15127 => std_logic_vector(to_unsigned( 48,8)),
			15128 => std_logic_vector(to_unsigned( 25,8)),
			15129 => std_logic_vector(to_unsigned( 136,8)),
			15130 => std_logic_vector(to_unsigned( 8,8)),
			15131 => std_logic_vector(to_unsigned( 230,8)),
			15132 => std_logic_vector(to_unsigned( 22,8)),
			15133 => std_logic_vector(to_unsigned( 3,8)),
			15134 => std_logic_vector(to_unsigned( 222,8)),
			15135 => std_logic_vector(to_unsigned( 77,8)),
			15136 => std_logic_vector(to_unsigned( 38,8)),
			15137 => std_logic_vector(to_unsigned( 53,8)),
			15138 => std_logic_vector(to_unsigned( 7,8)),
			15139 => std_logic_vector(to_unsigned( 206,8)),
			15140 => std_logic_vector(to_unsigned( 63,8)),
			15141 => std_logic_vector(to_unsigned( 65,8)),
			15142 => std_logic_vector(to_unsigned( 131,8)),
			15143 => std_logic_vector(to_unsigned( 186,8)),
			15144 => std_logic_vector(to_unsigned( 249,8)),
			15145 => std_logic_vector(to_unsigned( 12,8)),
			15146 => std_logic_vector(to_unsigned( 45,8)),
			15147 => std_logic_vector(to_unsigned( 196,8)),
			15148 => std_logic_vector(to_unsigned( 128,8)),
			15149 => std_logic_vector(to_unsigned( 33,8)),
			15150 => std_logic_vector(to_unsigned( 93,8)),
			15151 => std_logic_vector(to_unsigned( 154,8)),
			15152 => std_logic_vector(to_unsigned( 95,8)),
			15153 => std_logic_vector(to_unsigned( 126,8)),
			15154 => std_logic_vector(to_unsigned( 155,8)),
			15155 => std_logic_vector(to_unsigned( 99,8)),
			15156 => std_logic_vector(to_unsigned( 169,8)),
			15157 => std_logic_vector(to_unsigned( 44,8)),
			15158 => std_logic_vector(to_unsigned( 147,8)),
			15159 => std_logic_vector(to_unsigned( 192,8)),
			15160 => std_logic_vector(to_unsigned( 90,8)),
			15161 => std_logic_vector(to_unsigned( 19,8)),
			15162 => std_logic_vector(to_unsigned( 57,8)),
			15163 => std_logic_vector(to_unsigned( 85,8)),
			15164 => std_logic_vector(to_unsigned( 17,8)),
			15165 => std_logic_vector(to_unsigned( 134,8)),
			15166 => std_logic_vector(to_unsigned( 227,8)),
			15167 => std_logic_vector(to_unsigned( 0,8)),
			15168 => std_logic_vector(to_unsigned( 142,8)),
			15169 => std_logic_vector(to_unsigned( 96,8)),
			15170 => std_logic_vector(to_unsigned( 185,8)),
			15171 => std_logic_vector(to_unsigned( 118,8)),
			15172 => std_logic_vector(to_unsigned( 56,8)),
			15173 => std_logic_vector(to_unsigned( 12,8)),
			15174 => std_logic_vector(to_unsigned( 3,8)),
			15175 => std_logic_vector(to_unsigned( 43,8)),
			15176 => std_logic_vector(to_unsigned( 42,8)),
			15177 => std_logic_vector(to_unsigned( 253,8)),
			15178 => std_logic_vector(to_unsigned( 184,8)),
			15179 => std_logic_vector(to_unsigned( 51,8)),
			15180 => std_logic_vector(to_unsigned( 140,8)),
			15181 => std_logic_vector(to_unsigned( 176,8)),
			15182 => std_logic_vector(to_unsigned( 83,8)),
			15183 => std_logic_vector(to_unsigned( 19,8)),
			15184 => std_logic_vector(to_unsigned( 63,8)),
			15185 => std_logic_vector(to_unsigned( 254,8)),
			15186 => std_logic_vector(to_unsigned( 160,8)),
			15187 => std_logic_vector(to_unsigned( 244,8)),
			15188 => std_logic_vector(to_unsigned( 31,8)),
			15189 => std_logic_vector(to_unsigned( 95,8)),
			15190 => std_logic_vector(to_unsigned( 233,8)),
			15191 => std_logic_vector(to_unsigned( 182,8)),
			15192 => std_logic_vector(to_unsigned( 110,8)),
			15193 => std_logic_vector(to_unsigned( 240,8)),
			15194 => std_logic_vector(to_unsigned( 209,8)),
			15195 => std_logic_vector(to_unsigned( 53,8)),
			15196 => std_logic_vector(to_unsigned( 18,8)),
			15197 => std_logic_vector(to_unsigned( 245,8)),
			15198 => std_logic_vector(to_unsigned( 183,8)),
			15199 => std_logic_vector(to_unsigned( 113,8)),
			15200 => std_logic_vector(to_unsigned( 252,8)),
			15201 => std_logic_vector(to_unsigned( 179,8)),
			15202 => std_logic_vector(to_unsigned( 70,8)),
			15203 => std_logic_vector(to_unsigned( 61,8)),
			15204 => std_logic_vector(to_unsigned( 146,8)),
			15205 => std_logic_vector(to_unsigned( 125,8)),
			15206 => std_logic_vector(to_unsigned( 96,8)),
			15207 => std_logic_vector(to_unsigned( 55,8)),
			15208 => std_logic_vector(to_unsigned( 116,8)),
			15209 => std_logic_vector(to_unsigned( 89,8)),
			15210 => std_logic_vector(to_unsigned( 132,8)),
			15211 => std_logic_vector(to_unsigned( 158,8)),
			15212 => std_logic_vector(to_unsigned( 23,8)),
			15213 => std_logic_vector(to_unsigned( 255,8)),
			15214 => std_logic_vector(to_unsigned( 33,8)),
			15215 => std_logic_vector(to_unsigned( 55,8)),
			15216 => std_logic_vector(to_unsigned( 108,8)),
			15217 => std_logic_vector(to_unsigned( 37,8)),
			15218 => std_logic_vector(to_unsigned( 3,8)),
			15219 => std_logic_vector(to_unsigned( 33,8)),
			15220 => std_logic_vector(to_unsigned( 190,8)),
			15221 => std_logic_vector(to_unsigned( 189,8)),
			15222 => std_logic_vector(to_unsigned( 10,8)),
			15223 => std_logic_vector(to_unsigned( 114,8)),
			15224 => std_logic_vector(to_unsigned( 224,8)),
			15225 => std_logic_vector(to_unsigned( 134,8)),
			15226 => std_logic_vector(to_unsigned( 142,8)),
			15227 => std_logic_vector(to_unsigned( 17,8)),
			15228 => std_logic_vector(to_unsigned( 29,8)),
			15229 => std_logic_vector(to_unsigned( 227,8)),
			15230 => std_logic_vector(to_unsigned( 216,8)),
			15231 => std_logic_vector(to_unsigned( 249,8)),
			15232 => std_logic_vector(to_unsigned( 12,8)),
			15233 => std_logic_vector(to_unsigned( 169,8)),
			15234 => std_logic_vector(to_unsigned( 86,8)),
			15235 => std_logic_vector(to_unsigned( 127,8)),
			15236 => std_logic_vector(to_unsigned( 79,8)),
			15237 => std_logic_vector(to_unsigned( 244,8)),
			15238 => std_logic_vector(to_unsigned( 125,8)),
			15239 => std_logic_vector(to_unsigned( 127,8)),
			15240 => std_logic_vector(to_unsigned( 192,8)),
			15241 => std_logic_vector(to_unsigned( 124,8)),
			15242 => std_logic_vector(to_unsigned( 198,8)),
			15243 => std_logic_vector(to_unsigned( 64,8)),
			15244 => std_logic_vector(to_unsigned( 54,8)),
			15245 => std_logic_vector(to_unsigned( 234,8)),
			15246 => std_logic_vector(to_unsigned( 119,8)),
			15247 => std_logic_vector(to_unsigned( 122,8)),
			15248 => std_logic_vector(to_unsigned( 235,8)),
			15249 => std_logic_vector(to_unsigned( 217,8)),
			15250 => std_logic_vector(to_unsigned( 106,8)),
			15251 => std_logic_vector(to_unsigned( 88,8)),
			15252 => std_logic_vector(to_unsigned( 44,8)),
			15253 => std_logic_vector(to_unsigned( 167,8)),
			15254 => std_logic_vector(to_unsigned( 157,8)),
			15255 => std_logic_vector(to_unsigned( 18,8)),
			15256 => std_logic_vector(to_unsigned( 66,8)),
			15257 => std_logic_vector(to_unsigned( 175,8)),
			15258 => std_logic_vector(to_unsigned( 64,8)),
			15259 => std_logic_vector(to_unsigned( 65,8)),
			15260 => std_logic_vector(to_unsigned( 106,8)),
			15261 => std_logic_vector(to_unsigned( 158,8)),
			15262 => std_logic_vector(to_unsigned( 51,8)),
			15263 => std_logic_vector(to_unsigned( 243,8)),
			15264 => std_logic_vector(to_unsigned( 93,8)),
			15265 => std_logic_vector(to_unsigned( 70,8)),
			15266 => std_logic_vector(to_unsigned( 88,8)),
			15267 => std_logic_vector(to_unsigned( 58,8)),
			15268 => std_logic_vector(to_unsigned( 213,8)),
			15269 => std_logic_vector(to_unsigned( 2,8)),
			15270 => std_logic_vector(to_unsigned( 186,8)),
			15271 => std_logic_vector(to_unsigned( 37,8)),
			15272 => std_logic_vector(to_unsigned( 166,8)),
			15273 => std_logic_vector(to_unsigned( 175,8)),
			15274 => std_logic_vector(to_unsigned( 86,8)),
			15275 => std_logic_vector(to_unsigned( 130,8)),
			15276 => std_logic_vector(to_unsigned( 58,8)),
			15277 => std_logic_vector(to_unsigned( 203,8)),
			15278 => std_logic_vector(to_unsigned( 175,8)),
			15279 => std_logic_vector(to_unsigned( 76,8)),
			15280 => std_logic_vector(to_unsigned( 21,8)),
			15281 => std_logic_vector(to_unsigned( 128,8)),
			15282 => std_logic_vector(to_unsigned( 149,8)),
			15283 => std_logic_vector(to_unsigned( 130,8)),
			15284 => std_logic_vector(to_unsigned( 202,8)),
			15285 => std_logic_vector(to_unsigned( 240,8)),
			15286 => std_logic_vector(to_unsigned( 32,8)),
			15287 => std_logic_vector(to_unsigned( 234,8)),
			15288 => std_logic_vector(to_unsigned( 173,8)),
			15289 => std_logic_vector(to_unsigned( 147,8)),
			15290 => std_logic_vector(to_unsigned( 186,8)),
			15291 => std_logic_vector(to_unsigned( 2,8)),
			15292 => std_logic_vector(to_unsigned( 224,8)),
			15293 => std_logic_vector(to_unsigned( 106,8)),
			15294 => std_logic_vector(to_unsigned( 28,8)),
			15295 => std_logic_vector(to_unsigned( 148,8)),
			15296 => std_logic_vector(to_unsigned( 218,8)),
			15297 => std_logic_vector(to_unsigned( 73,8)),
			15298 => std_logic_vector(to_unsigned( 122,8)),
			15299 => std_logic_vector(to_unsigned( 56,8)),
			15300 => std_logic_vector(to_unsigned( 80,8)),
			15301 => std_logic_vector(to_unsigned( 83,8)),
			15302 => std_logic_vector(to_unsigned( 116,8)),
			15303 => std_logic_vector(to_unsigned( 0,8)),
			15304 => std_logic_vector(to_unsigned( 2,8)),
			15305 => std_logic_vector(to_unsigned( 155,8)),
			15306 => std_logic_vector(to_unsigned( 153,8)),
			15307 => std_logic_vector(to_unsigned( 205,8)),
			15308 => std_logic_vector(to_unsigned( 182,8)),
			15309 => std_logic_vector(to_unsigned( 179,8)),
			15310 => std_logic_vector(to_unsigned( 129,8)),
			15311 => std_logic_vector(to_unsigned( 225,8)),
			15312 => std_logic_vector(to_unsigned( 48,8)),
			15313 => std_logic_vector(to_unsigned( 203,8)),
			15314 => std_logic_vector(to_unsigned( 35,8)),
			15315 => std_logic_vector(to_unsigned( 247,8)),
			15316 => std_logic_vector(to_unsigned( 78,8)),
			15317 => std_logic_vector(to_unsigned( 20,8)),
			15318 => std_logic_vector(to_unsigned( 74,8)),
			15319 => std_logic_vector(to_unsigned( 5,8)),
			15320 => std_logic_vector(to_unsigned( 6,8)),
			15321 => std_logic_vector(to_unsigned( 152,8)),
			15322 => std_logic_vector(to_unsigned( 137,8)),
			15323 => std_logic_vector(to_unsigned( 219,8)),
			15324 => std_logic_vector(to_unsigned( 46,8)),
			15325 => std_logic_vector(to_unsigned( 227,8)),
			15326 => std_logic_vector(to_unsigned( 194,8)),
			15327 => std_logic_vector(to_unsigned( 213,8)),
			15328 => std_logic_vector(to_unsigned( 241,8)),
			15329 => std_logic_vector(to_unsigned( 26,8)),
			15330 => std_logic_vector(to_unsigned( 38,8)),
			15331 => std_logic_vector(to_unsigned( 2,8)),
			15332 => std_logic_vector(to_unsigned( 136,8)),
			15333 => std_logic_vector(to_unsigned( 185,8)),
			15334 => std_logic_vector(to_unsigned( 66,8)),
			15335 => std_logic_vector(to_unsigned( 15,8)),
			15336 => std_logic_vector(to_unsigned( 255,8)),
			15337 => std_logic_vector(to_unsigned( 252,8)),
			15338 => std_logic_vector(to_unsigned( 99,8)),
			15339 => std_logic_vector(to_unsigned( 34,8)),
			15340 => std_logic_vector(to_unsigned( 76,8)),
			15341 => std_logic_vector(to_unsigned( 83,8)),
			15342 => std_logic_vector(to_unsigned( 1,8)),
			15343 => std_logic_vector(to_unsigned( 75,8)),
			15344 => std_logic_vector(to_unsigned( 80,8)),
			15345 => std_logic_vector(to_unsigned( 70,8)),
			15346 => std_logic_vector(to_unsigned( 151,8)),
			15347 => std_logic_vector(to_unsigned( 71,8)),
			15348 => std_logic_vector(to_unsigned( 68,8)),
			15349 => std_logic_vector(to_unsigned( 209,8)),
			15350 => std_logic_vector(to_unsigned( 12,8)),
			15351 => std_logic_vector(to_unsigned( 233,8)),
			15352 => std_logic_vector(to_unsigned( 229,8)),
			15353 => std_logic_vector(to_unsigned( 6,8)),
			15354 => std_logic_vector(to_unsigned( 208,8)),
			15355 => std_logic_vector(to_unsigned( 240,8)),
			15356 => std_logic_vector(to_unsigned( 245,8)),
			15357 => std_logic_vector(to_unsigned( 43,8)),
			15358 => std_logic_vector(to_unsigned( 95,8)),
			15359 => std_logic_vector(to_unsigned( 26,8)),
			15360 => std_logic_vector(to_unsigned( 121,8)),
			15361 => std_logic_vector(to_unsigned( 143,8)),
			15362 => std_logic_vector(to_unsigned( 205,8)),
			15363 => std_logic_vector(to_unsigned( 181,8)),
			15364 => std_logic_vector(to_unsigned( 198,8)),
			15365 => std_logic_vector(to_unsigned( 236,8)),
			15366 => std_logic_vector(to_unsigned( 134,8)),
			15367 => std_logic_vector(to_unsigned( 130,8)),
			15368 => std_logic_vector(to_unsigned( 40,8)),
			15369 => std_logic_vector(to_unsigned( 26,8)),
			15370 => std_logic_vector(to_unsigned( 94,8)),
			15371 => std_logic_vector(to_unsigned( 167,8)),
			15372 => std_logic_vector(to_unsigned( 146,8)),
			15373 => std_logic_vector(to_unsigned( 74,8)),
			15374 => std_logic_vector(to_unsigned( 28,8)),
			15375 => std_logic_vector(to_unsigned( 4,8)),
			15376 => std_logic_vector(to_unsigned( 101,8)),
			15377 => std_logic_vector(to_unsigned( 63,8)),
			15378 => std_logic_vector(to_unsigned( 6,8)),
			15379 => std_logic_vector(to_unsigned( 17,8)),
			15380 => std_logic_vector(to_unsigned( 208,8)),
			15381 => std_logic_vector(to_unsigned( 108,8)),
			15382 => std_logic_vector(to_unsigned( 183,8)),
			15383 => std_logic_vector(to_unsigned( 101,8)),
			15384 => std_logic_vector(to_unsigned( 10,8)),
			15385 => std_logic_vector(to_unsigned( 60,8)),
			15386 => std_logic_vector(to_unsigned( 139,8)),
			15387 => std_logic_vector(to_unsigned( 78,8)),
			15388 => std_logic_vector(to_unsigned( 135,8)),
			15389 => std_logic_vector(to_unsigned( 221,8)),
			15390 => std_logic_vector(to_unsigned( 58,8)),
			15391 => std_logic_vector(to_unsigned( 131,8)),
			15392 => std_logic_vector(to_unsigned( 172,8)),
			15393 => std_logic_vector(to_unsigned( 178,8)),
			15394 => std_logic_vector(to_unsigned( 123,8)),
			15395 => std_logic_vector(to_unsigned( 112,8)),
			15396 => std_logic_vector(to_unsigned( 156,8)),
			15397 => std_logic_vector(to_unsigned( 151,8)),
			15398 => std_logic_vector(to_unsigned( 66,8)),
			15399 => std_logic_vector(to_unsigned( 163,8)),
			15400 => std_logic_vector(to_unsigned( 6,8)),
			15401 => std_logic_vector(to_unsigned( 238,8)),
			15402 => std_logic_vector(to_unsigned( 136,8)),
			15403 => std_logic_vector(to_unsigned( 164,8)),
			15404 => std_logic_vector(to_unsigned( 153,8)),
			15405 => std_logic_vector(to_unsigned( 162,8)),
			15406 => std_logic_vector(to_unsigned( 176,8)),
			15407 => std_logic_vector(to_unsigned( 186,8)),
			15408 => std_logic_vector(to_unsigned( 12,8)),
			15409 => std_logic_vector(to_unsigned( 138,8)),
			15410 => std_logic_vector(to_unsigned( 231,8)),
			15411 => std_logic_vector(to_unsigned( 177,8)),
			15412 => std_logic_vector(to_unsigned( 220,8)),
			15413 => std_logic_vector(to_unsigned( 4,8)),
			15414 => std_logic_vector(to_unsigned( 227,8)),
			15415 => std_logic_vector(to_unsigned( 126,8)),
			15416 => std_logic_vector(to_unsigned( 189,8)),
			15417 => std_logic_vector(to_unsigned( 157,8)),
			15418 => std_logic_vector(to_unsigned( 12,8)),
			15419 => std_logic_vector(to_unsigned( 202,8)),
			15420 => std_logic_vector(to_unsigned( 104,8)),
			15421 => std_logic_vector(to_unsigned( 99,8)),
			15422 => std_logic_vector(to_unsigned( 216,8)),
			15423 => std_logic_vector(to_unsigned( 153,8)),
			15424 => std_logic_vector(to_unsigned( 25,8)),
			15425 => std_logic_vector(to_unsigned( 49,8)),
			15426 => std_logic_vector(to_unsigned( 86,8)),
			15427 => std_logic_vector(to_unsigned( 208,8)),
			15428 => std_logic_vector(to_unsigned( 217,8)),
			15429 => std_logic_vector(to_unsigned( 104,8)),
			15430 => std_logic_vector(to_unsigned( 140,8)),
			15431 => std_logic_vector(to_unsigned( 226,8)),
			15432 => std_logic_vector(to_unsigned( 32,8)),
			15433 => std_logic_vector(to_unsigned( 8,8)),
			15434 => std_logic_vector(to_unsigned( 36,8)),
			15435 => std_logic_vector(to_unsigned( 66,8)),
			15436 => std_logic_vector(to_unsigned( 38,8)),
			15437 => std_logic_vector(to_unsigned( 40,8)),
			15438 => std_logic_vector(to_unsigned( 159,8)),
			15439 => std_logic_vector(to_unsigned( 123,8)),
			15440 => std_logic_vector(to_unsigned( 72,8)),
			15441 => std_logic_vector(to_unsigned( 153,8)),
			15442 => std_logic_vector(to_unsigned( 156,8)),
			15443 => std_logic_vector(to_unsigned( 47,8)),
			15444 => std_logic_vector(to_unsigned( 199,8)),
			15445 => std_logic_vector(to_unsigned( 244,8)),
			15446 => std_logic_vector(to_unsigned( 86,8)),
			15447 => std_logic_vector(to_unsigned( 227,8)),
			15448 => std_logic_vector(to_unsigned( 24,8)),
			15449 => std_logic_vector(to_unsigned( 186,8)),
			15450 => std_logic_vector(to_unsigned( 208,8)),
			15451 => std_logic_vector(to_unsigned( 61,8)),
			15452 => std_logic_vector(to_unsigned( 162,8)),
			15453 => std_logic_vector(to_unsigned( 185,8)),
			15454 => std_logic_vector(to_unsigned( 203,8)),
			15455 => std_logic_vector(to_unsigned( 116,8)),
			15456 => std_logic_vector(to_unsigned( 199,8)),
			15457 => std_logic_vector(to_unsigned( 102,8)),
			15458 => std_logic_vector(to_unsigned( 169,8)),
			15459 => std_logic_vector(to_unsigned( 137,8)),
			15460 => std_logic_vector(to_unsigned( 138,8)),
			15461 => std_logic_vector(to_unsigned( 52,8)),
			15462 => std_logic_vector(to_unsigned( 133,8)),
			15463 => std_logic_vector(to_unsigned( 66,8)),
			15464 => std_logic_vector(to_unsigned( 175,8)),
			15465 => std_logic_vector(to_unsigned( 115,8)),
			15466 => std_logic_vector(to_unsigned( 8,8)),
			15467 => std_logic_vector(to_unsigned( 254,8)),
			15468 => std_logic_vector(to_unsigned( 173,8)),
			15469 => std_logic_vector(to_unsigned( 163,8)),
			15470 => std_logic_vector(to_unsigned( 22,8)),
			15471 => std_logic_vector(to_unsigned( 52,8)),
			15472 => std_logic_vector(to_unsigned( 49,8)),
			15473 => std_logic_vector(to_unsigned( 168,8)),
			15474 => std_logic_vector(to_unsigned( 247,8)),
			15475 => std_logic_vector(to_unsigned( 207,8)),
			15476 => std_logic_vector(to_unsigned( 193,8)),
			15477 => std_logic_vector(to_unsigned( 67,8)),
			15478 => std_logic_vector(to_unsigned( 194,8)),
			15479 => std_logic_vector(to_unsigned( 101,8)),
			15480 => std_logic_vector(to_unsigned( 40,8)),
			15481 => std_logic_vector(to_unsigned( 168,8)),
			15482 => std_logic_vector(to_unsigned( 35,8)),
			15483 => std_logic_vector(to_unsigned( 8,8)),
			15484 => std_logic_vector(to_unsigned( 224,8)),
			15485 => std_logic_vector(to_unsigned( 152,8)),
			15486 => std_logic_vector(to_unsigned( 180,8)),
			15487 => std_logic_vector(to_unsigned( 202,8)),
			15488 => std_logic_vector(to_unsigned( 18,8)),
			15489 => std_logic_vector(to_unsigned( 140,8)),
			15490 => std_logic_vector(to_unsigned( 194,8)),
			15491 => std_logic_vector(to_unsigned( 202,8)),
			15492 => std_logic_vector(to_unsigned( 222,8)),
			15493 => std_logic_vector(to_unsigned( 214,8)),
			15494 => std_logic_vector(to_unsigned( 240,8)),
			15495 => std_logic_vector(to_unsigned( 149,8)),
			15496 => std_logic_vector(to_unsigned( 231,8)),
			15497 => std_logic_vector(to_unsigned( 140,8)),
			15498 => std_logic_vector(to_unsigned( 27,8)),
			15499 => std_logic_vector(to_unsigned( 96,8)),
			15500 => std_logic_vector(to_unsigned( 228,8)),
			15501 => std_logic_vector(to_unsigned( 107,8)),
			15502 => std_logic_vector(to_unsigned( 237,8)),
			15503 => std_logic_vector(to_unsigned( 112,8)),
			15504 => std_logic_vector(to_unsigned( 179,8)),
			15505 => std_logic_vector(to_unsigned( 0,8)),
			15506 => std_logic_vector(to_unsigned( 197,8)),
			15507 => std_logic_vector(to_unsigned( 178,8)),
			15508 => std_logic_vector(to_unsigned( 122,8)),
			15509 => std_logic_vector(to_unsigned( 18,8)),
			15510 => std_logic_vector(to_unsigned( 107,8)),
			15511 => std_logic_vector(to_unsigned( 205,8)),
			15512 => std_logic_vector(to_unsigned( 224,8)),
			15513 => std_logic_vector(to_unsigned( 176,8)),
			15514 => std_logic_vector(to_unsigned( 118,8)),
			15515 => std_logic_vector(to_unsigned( 253,8)),
			15516 => std_logic_vector(to_unsigned( 43,8)),
			15517 => std_logic_vector(to_unsigned( 3,8)),
			15518 => std_logic_vector(to_unsigned( 133,8)),
			15519 => std_logic_vector(to_unsigned( 100,8)),
			15520 => std_logic_vector(to_unsigned( 113,8)),
			15521 => std_logic_vector(to_unsigned( 16,8)),
			15522 => std_logic_vector(to_unsigned( 184,8)),
			15523 => std_logic_vector(to_unsigned( 119,8)),
			15524 => std_logic_vector(to_unsigned( 63,8)),
			15525 => std_logic_vector(to_unsigned( 200,8)),
			15526 => std_logic_vector(to_unsigned( 231,8)),
			15527 => std_logic_vector(to_unsigned( 140,8)),
			15528 => std_logic_vector(to_unsigned( 92,8)),
			15529 => std_logic_vector(to_unsigned( 116,8)),
			15530 => std_logic_vector(to_unsigned( 171,8)),
			15531 => std_logic_vector(to_unsigned( 89,8)),
			15532 => std_logic_vector(to_unsigned( 177,8)),
			15533 => std_logic_vector(to_unsigned( 18,8)),
			15534 => std_logic_vector(to_unsigned( 22,8)),
			15535 => std_logic_vector(to_unsigned( 39,8)),
			15536 => std_logic_vector(to_unsigned( 196,8)),
			15537 => std_logic_vector(to_unsigned( 155,8)),
			15538 => std_logic_vector(to_unsigned( 189,8)),
			15539 => std_logic_vector(to_unsigned( 75,8)),
			15540 => std_logic_vector(to_unsigned( 216,8)),
			15541 => std_logic_vector(to_unsigned( 192,8)),
			15542 => std_logic_vector(to_unsigned( 218,8)),
			15543 => std_logic_vector(to_unsigned( 69,8)),
			15544 => std_logic_vector(to_unsigned( 58,8)),
			15545 => std_logic_vector(to_unsigned( 155,8)),
			15546 => std_logic_vector(to_unsigned( 223,8)),
			15547 => std_logic_vector(to_unsigned( 189,8)),
			15548 => std_logic_vector(to_unsigned( 63,8)),
			15549 => std_logic_vector(to_unsigned( 17,8)),
			15550 => std_logic_vector(to_unsigned( 116,8)),
			15551 => std_logic_vector(to_unsigned( 54,8)),
			15552 => std_logic_vector(to_unsigned( 104,8)),
			15553 => std_logic_vector(to_unsigned( 10,8)),
			15554 => std_logic_vector(to_unsigned( 196,8)),
			15555 => std_logic_vector(to_unsigned( 66,8)),
			15556 => std_logic_vector(to_unsigned( 212,8)),
			15557 => std_logic_vector(to_unsigned( 158,8)),
			15558 => std_logic_vector(to_unsigned( 89,8)),
			15559 => std_logic_vector(to_unsigned( 189,8)),
			15560 => std_logic_vector(to_unsigned( 210,8)),
			15561 => std_logic_vector(to_unsigned( 125,8)),
			15562 => std_logic_vector(to_unsigned( 158,8)),
			15563 => std_logic_vector(to_unsigned( 166,8)),
			15564 => std_logic_vector(to_unsigned( 232,8)),
			15565 => std_logic_vector(to_unsigned( 244,8)),
			15566 => std_logic_vector(to_unsigned( 82,8)),
			15567 => std_logic_vector(to_unsigned( 234,8)),
			15568 => std_logic_vector(to_unsigned( 127,8)),
			15569 => std_logic_vector(to_unsigned( 141,8)),
			15570 => std_logic_vector(to_unsigned( 53,8)),
			15571 => std_logic_vector(to_unsigned( 33,8)),
			15572 => std_logic_vector(to_unsigned( 34,8)),
			15573 => std_logic_vector(to_unsigned( 226,8)),
			15574 => std_logic_vector(to_unsigned( 44,8)),
			15575 => std_logic_vector(to_unsigned( 61,8)),
			15576 => std_logic_vector(to_unsigned( 252,8)),
			15577 => std_logic_vector(to_unsigned( 83,8)),
			15578 => std_logic_vector(to_unsigned( 126,8)),
			15579 => std_logic_vector(to_unsigned( 193,8)),
			15580 => std_logic_vector(to_unsigned( 139,8)),
			15581 => std_logic_vector(to_unsigned( 207,8)),
			15582 => std_logic_vector(to_unsigned( 118,8)),
			15583 => std_logic_vector(to_unsigned( 47,8)),
			15584 => std_logic_vector(to_unsigned( 205,8)),
			15585 => std_logic_vector(to_unsigned( 3,8)),
			15586 => std_logic_vector(to_unsigned( 226,8)),
			15587 => std_logic_vector(to_unsigned( 88,8)),
			15588 => std_logic_vector(to_unsigned( 211,8)),
			15589 => std_logic_vector(to_unsigned( 19,8)),
			15590 => std_logic_vector(to_unsigned( 187,8)),
			15591 => std_logic_vector(to_unsigned( 143,8)),
			15592 => std_logic_vector(to_unsigned( 25,8)),
			15593 => std_logic_vector(to_unsigned( 175,8)),
			15594 => std_logic_vector(to_unsigned( 16,8)),
			15595 => std_logic_vector(to_unsigned( 12,8)),
			15596 => std_logic_vector(to_unsigned( 140,8)),
			15597 => std_logic_vector(to_unsigned( 28,8)),
			15598 => std_logic_vector(to_unsigned( 104,8)),
			15599 => std_logic_vector(to_unsigned( 69,8)),
			15600 => std_logic_vector(to_unsigned( 250,8)),
			15601 => std_logic_vector(to_unsigned( 21,8)),
			15602 => std_logic_vector(to_unsigned( 16,8)),
			15603 => std_logic_vector(to_unsigned( 35,8)),
			15604 => std_logic_vector(to_unsigned( 81,8)),
			15605 => std_logic_vector(to_unsigned( 94,8)),
			15606 => std_logic_vector(to_unsigned( 103,8)),
			15607 => std_logic_vector(to_unsigned( 162,8)),
			15608 => std_logic_vector(to_unsigned( 229,8)),
			15609 => std_logic_vector(to_unsigned( 238,8)),
			15610 => std_logic_vector(to_unsigned( 93,8)),
			15611 => std_logic_vector(to_unsigned( 180,8)),
			15612 => std_logic_vector(to_unsigned( 243,8)),
			15613 => std_logic_vector(to_unsigned( 164,8)),
			15614 => std_logic_vector(to_unsigned( 57,8)),
			15615 => std_logic_vector(to_unsigned( 165,8)),
			15616 => std_logic_vector(to_unsigned( 203,8)),
			15617 => std_logic_vector(to_unsigned( 239,8)),
			15618 => std_logic_vector(to_unsigned( 201,8)),
			15619 => std_logic_vector(to_unsigned( 142,8)),
			15620 => std_logic_vector(to_unsigned( 175,8)),
			15621 => std_logic_vector(to_unsigned( 217,8)),
			15622 => std_logic_vector(to_unsigned( 50,8)),
			15623 => std_logic_vector(to_unsigned( 89,8)),
			15624 => std_logic_vector(to_unsigned( 113,8)),
			15625 => std_logic_vector(to_unsigned( 240,8)),
			15626 => std_logic_vector(to_unsigned( 169,8)),
			15627 => std_logic_vector(to_unsigned( 246,8)),
			15628 => std_logic_vector(to_unsigned( 188,8)),
			15629 => std_logic_vector(to_unsigned( 1,8)),
			15630 => std_logic_vector(to_unsigned( 165,8)),
			15631 => std_logic_vector(to_unsigned( 100,8)),
			15632 => std_logic_vector(to_unsigned( 30,8)),
			15633 => std_logic_vector(to_unsigned( 228,8)),
			15634 => std_logic_vector(to_unsigned( 135,8)),
			15635 => std_logic_vector(to_unsigned( 243,8)),
			15636 => std_logic_vector(to_unsigned( 147,8)),
			15637 => std_logic_vector(to_unsigned( 189,8)),
			15638 => std_logic_vector(to_unsigned( 238,8)),
			15639 => std_logic_vector(to_unsigned( 64,8)),
			15640 => std_logic_vector(to_unsigned( 36,8)),
			15641 => std_logic_vector(to_unsigned( 115,8)),
			15642 => std_logic_vector(to_unsigned( 9,8)),
			15643 => std_logic_vector(to_unsigned( 115,8)),
			15644 => std_logic_vector(to_unsigned( 174,8)),
			15645 => std_logic_vector(to_unsigned( 36,8)),
			15646 => std_logic_vector(to_unsigned( 84,8)),
			15647 => std_logic_vector(to_unsigned( 208,8)),
			15648 => std_logic_vector(to_unsigned( 248,8)),
			15649 => std_logic_vector(to_unsigned( 51,8)),
			15650 => std_logic_vector(to_unsigned( 106,8)),
			15651 => std_logic_vector(to_unsigned( 47,8)),
			15652 => std_logic_vector(to_unsigned( 136,8)),
			15653 => std_logic_vector(to_unsigned( 78,8)),
			15654 => std_logic_vector(to_unsigned( 42,8)),
			15655 => std_logic_vector(to_unsigned( 183,8)),
			15656 => std_logic_vector(to_unsigned( 183,8)),
			15657 => std_logic_vector(to_unsigned( 125,8)),
			15658 => std_logic_vector(to_unsigned( 187,8)),
			15659 => std_logic_vector(to_unsigned( 22,8)),
			15660 => std_logic_vector(to_unsigned( 230,8)),
			15661 => std_logic_vector(to_unsigned( 106,8)),
			15662 => std_logic_vector(to_unsigned( 81,8)),
			15663 => std_logic_vector(to_unsigned( 205,8)),
			15664 => std_logic_vector(to_unsigned( 12,8)),
			15665 => std_logic_vector(to_unsigned( 22,8)),
			15666 => std_logic_vector(to_unsigned( 9,8)),
			15667 => std_logic_vector(to_unsigned( 137,8)),
			15668 => std_logic_vector(to_unsigned( 159,8)),
			15669 => std_logic_vector(to_unsigned( 16,8)),
			15670 => std_logic_vector(to_unsigned( 137,8)),
			15671 => std_logic_vector(to_unsigned( 252,8)),
			15672 => std_logic_vector(to_unsigned( 150,8)),
			15673 => std_logic_vector(to_unsigned( 161,8)),
			15674 => std_logic_vector(to_unsigned( 87,8)),
			15675 => std_logic_vector(to_unsigned( 124,8)),
			15676 => std_logic_vector(to_unsigned( 183,8)),
			15677 => std_logic_vector(to_unsigned( 236,8)),
			15678 => std_logic_vector(to_unsigned( 113,8)),
			15679 => std_logic_vector(to_unsigned( 8,8)),
			15680 => std_logic_vector(to_unsigned( 242,8)),
			15681 => std_logic_vector(to_unsigned( 77,8)),
			15682 => std_logic_vector(to_unsigned( 42,8)),
			15683 => std_logic_vector(to_unsigned( 146,8)),
			15684 => std_logic_vector(to_unsigned( 134,8)),
			15685 => std_logic_vector(to_unsigned( 167,8)),
			15686 => std_logic_vector(to_unsigned( 123,8)),
			15687 => std_logic_vector(to_unsigned( 230,8)),
			15688 => std_logic_vector(to_unsigned( 185,8)),
			15689 => std_logic_vector(to_unsigned( 223,8)),
			15690 => std_logic_vector(to_unsigned( 12,8)),
			15691 => std_logic_vector(to_unsigned( 70,8)),
			15692 => std_logic_vector(to_unsigned( 108,8)),
			15693 => std_logic_vector(to_unsigned( 253,8)),
			15694 => std_logic_vector(to_unsigned( 202,8)),
			15695 => std_logic_vector(to_unsigned( 117,8)),
			15696 => std_logic_vector(to_unsigned( 62,8)),
			15697 => std_logic_vector(to_unsigned( 161,8)),
			15698 => std_logic_vector(to_unsigned( 208,8)),
			15699 => std_logic_vector(to_unsigned( 201,8)),
			15700 => std_logic_vector(to_unsigned( 71,8)),
			15701 => std_logic_vector(to_unsigned( 177,8)),
			15702 => std_logic_vector(to_unsigned( 159,8)),
			15703 => std_logic_vector(to_unsigned( 55,8)),
			15704 => std_logic_vector(to_unsigned( 76,8)),
			15705 => std_logic_vector(to_unsigned( 169,8)),
			15706 => std_logic_vector(to_unsigned( 142,8)),
			15707 => std_logic_vector(to_unsigned( 119,8)),
			15708 => std_logic_vector(to_unsigned( 68,8)),
			15709 => std_logic_vector(to_unsigned( 31,8)),
			15710 => std_logic_vector(to_unsigned( 23,8)),
			15711 => std_logic_vector(to_unsigned( 150,8)),
			15712 => std_logic_vector(to_unsigned( 30,8)),
			15713 => std_logic_vector(to_unsigned( 125,8)),
			15714 => std_logic_vector(to_unsigned( 189,8)),
			15715 => std_logic_vector(to_unsigned( 209,8)),
			15716 => std_logic_vector(to_unsigned( 132,8)),
			15717 => std_logic_vector(to_unsigned( 182,8)),
			15718 => std_logic_vector(to_unsigned( 201,8)),
			15719 => std_logic_vector(to_unsigned( 129,8)),
			15720 => std_logic_vector(to_unsigned( 224,8)),
			15721 => std_logic_vector(to_unsigned( 1,8)),
			15722 => std_logic_vector(to_unsigned( 102,8)),
			15723 => std_logic_vector(to_unsigned( 46,8)),
			15724 => std_logic_vector(to_unsigned( 180,8)),
			15725 => std_logic_vector(to_unsigned( 233,8)),
			15726 => std_logic_vector(to_unsigned( 147,8)),
			15727 => std_logic_vector(to_unsigned( 175,8)),
			15728 => std_logic_vector(to_unsigned( 94,8)),
			15729 => std_logic_vector(to_unsigned( 248,8)),
			15730 => std_logic_vector(to_unsigned( 197,8)),
			15731 => std_logic_vector(to_unsigned( 26,8)),
			15732 => std_logic_vector(to_unsigned( 84,8)),
			15733 => std_logic_vector(to_unsigned( 123,8)),
			15734 => std_logic_vector(to_unsigned( 126,8)),
			15735 => std_logic_vector(to_unsigned( 156,8)),
			15736 => std_logic_vector(to_unsigned( 249,8)),
			15737 => std_logic_vector(to_unsigned( 220,8)),
			15738 => std_logic_vector(to_unsigned( 57,8)),
			15739 => std_logic_vector(to_unsigned( 100,8)),
			15740 => std_logic_vector(to_unsigned( 32,8)),
			15741 => std_logic_vector(to_unsigned( 25,8)),
			15742 => std_logic_vector(to_unsigned( 38,8)),
			15743 => std_logic_vector(to_unsigned( 162,8)),
			15744 => std_logic_vector(to_unsigned( 253,8)),
			15745 => std_logic_vector(to_unsigned( 116,8)),
			15746 => std_logic_vector(to_unsigned( 68,8)),
			15747 => std_logic_vector(to_unsigned( 166,8)),
			15748 => std_logic_vector(to_unsigned( 202,8)),
			15749 => std_logic_vector(to_unsigned( 54,8)),
			15750 => std_logic_vector(to_unsigned( 8,8)),
			15751 => std_logic_vector(to_unsigned( 187,8)),
			15752 => std_logic_vector(to_unsigned( 76,8)),
			15753 => std_logic_vector(to_unsigned( 249,8)),
			15754 => std_logic_vector(to_unsigned( 25,8)),
			15755 => std_logic_vector(to_unsigned( 115,8)),
			15756 => std_logic_vector(to_unsigned( 27,8)),
			15757 => std_logic_vector(to_unsigned( 58,8)),
			15758 => std_logic_vector(to_unsigned( 200,8)),
			15759 => std_logic_vector(to_unsigned( 119,8)),
			15760 => std_logic_vector(to_unsigned( 25,8)),
			15761 => std_logic_vector(to_unsigned( 135,8)),
			15762 => std_logic_vector(to_unsigned( 219,8)),
			15763 => std_logic_vector(to_unsigned( 125,8)),
			15764 => std_logic_vector(to_unsigned( 107,8)),
			15765 => std_logic_vector(to_unsigned( 151,8)),
			15766 => std_logic_vector(to_unsigned( 104,8)),
			15767 => std_logic_vector(to_unsigned( 39,8)),
			15768 => std_logic_vector(to_unsigned( 15,8)),
			15769 => std_logic_vector(to_unsigned( 167,8)),
			15770 => std_logic_vector(to_unsigned( 95,8)),
			15771 => std_logic_vector(to_unsigned( 199,8)),
			15772 => std_logic_vector(to_unsigned( 225,8)),
			15773 => std_logic_vector(to_unsigned( 14,8)),
			15774 => std_logic_vector(to_unsigned( 96,8)),
			15775 => std_logic_vector(to_unsigned( 234,8)),
			15776 => std_logic_vector(to_unsigned( 223,8)),
			15777 => std_logic_vector(to_unsigned( 41,8)),
			15778 => std_logic_vector(to_unsigned( 234,8)),
			15779 => std_logic_vector(to_unsigned( 190,8)),
			15780 => std_logic_vector(to_unsigned( 117,8)),
			15781 => std_logic_vector(to_unsigned( 36,8)),
			15782 => std_logic_vector(to_unsigned( 164,8)),
			15783 => std_logic_vector(to_unsigned( 1,8)),
			15784 => std_logic_vector(to_unsigned( 19,8)),
			15785 => std_logic_vector(to_unsigned( 100,8)),
			15786 => std_logic_vector(to_unsigned( 23,8)),
			15787 => std_logic_vector(to_unsigned( 144,8)),
			15788 => std_logic_vector(to_unsigned( 84,8)),
			15789 => std_logic_vector(to_unsigned( 193,8)),
			15790 => std_logic_vector(to_unsigned( 110,8)),
			15791 => std_logic_vector(to_unsigned( 16,8)),
			15792 => std_logic_vector(to_unsigned( 187,8)),
			15793 => std_logic_vector(to_unsigned( 1,8)),
			15794 => std_logic_vector(to_unsigned( 191,8)),
			15795 => std_logic_vector(to_unsigned( 50,8)),
			15796 => std_logic_vector(to_unsigned( 124,8)),
			15797 => std_logic_vector(to_unsigned( 19,8)),
			15798 => std_logic_vector(to_unsigned( 217,8)),
			15799 => std_logic_vector(to_unsigned( 80,8)),
			15800 => std_logic_vector(to_unsigned( 19,8)),
			15801 => std_logic_vector(to_unsigned( 111,8)),
			15802 => std_logic_vector(to_unsigned( 179,8)),
			15803 => std_logic_vector(to_unsigned( 63,8)),
			15804 => std_logic_vector(to_unsigned( 113,8)),
			15805 => std_logic_vector(to_unsigned( 31,8)),
			15806 => std_logic_vector(to_unsigned( 4,8)),
			15807 => std_logic_vector(to_unsigned( 65,8)),
			15808 => std_logic_vector(to_unsigned( 0,8)),
			15809 => std_logic_vector(to_unsigned( 180,8)),
			15810 => std_logic_vector(to_unsigned( 131,8)),
			15811 => std_logic_vector(to_unsigned( 165,8)),
			15812 => std_logic_vector(to_unsigned( 219,8)),
			15813 => std_logic_vector(to_unsigned( 47,8)),
			15814 => std_logic_vector(to_unsigned( 134,8)),
			15815 => std_logic_vector(to_unsigned( 229,8)),
			15816 => std_logic_vector(to_unsigned( 252,8)),
			15817 => std_logic_vector(to_unsigned( 70,8)),
			15818 => std_logic_vector(to_unsigned( 176,8)),
			15819 => std_logic_vector(to_unsigned( 196,8)),
			15820 => std_logic_vector(to_unsigned( 237,8)),
			15821 => std_logic_vector(to_unsigned( 177,8)),
			15822 => std_logic_vector(to_unsigned( 59,8)),
			15823 => std_logic_vector(to_unsigned( 177,8)),
			15824 => std_logic_vector(to_unsigned( 110,8)),
			15825 => std_logic_vector(to_unsigned( 135,8)),
			15826 => std_logic_vector(to_unsigned( 251,8)),
			15827 => std_logic_vector(to_unsigned( 91,8)),
			15828 => std_logic_vector(to_unsigned( 188,8)),
			15829 => std_logic_vector(to_unsigned( 13,8)),
			15830 => std_logic_vector(to_unsigned( 191,8)),
			15831 => std_logic_vector(to_unsigned( 112,8)),
			15832 => std_logic_vector(to_unsigned( 84,8)),
			15833 => std_logic_vector(to_unsigned( 237,8)),
			15834 => std_logic_vector(to_unsigned( 12,8)),
			15835 => std_logic_vector(to_unsigned( 36,8)),
			15836 => std_logic_vector(to_unsigned( 44,8)),
			15837 => std_logic_vector(to_unsigned( 223,8)),
			15838 => std_logic_vector(to_unsigned( 58,8)),
			15839 => std_logic_vector(to_unsigned( 87,8)),
			15840 => std_logic_vector(to_unsigned( 218,8)),
			15841 => std_logic_vector(to_unsigned( 212,8)),
			15842 => std_logic_vector(to_unsigned( 96,8)),
			15843 => std_logic_vector(to_unsigned( 42,8)),
			15844 => std_logic_vector(to_unsigned( 40,8)),
			15845 => std_logic_vector(to_unsigned( 171,8)),
			15846 => std_logic_vector(to_unsigned( 225,8)),
			15847 => std_logic_vector(to_unsigned( 29,8)),
			15848 => std_logic_vector(to_unsigned( 133,8)),
			15849 => std_logic_vector(to_unsigned( 35,8)),
			15850 => std_logic_vector(to_unsigned( 90,8)),
			15851 => std_logic_vector(to_unsigned( 118,8)),
			15852 => std_logic_vector(to_unsigned( 46,8)),
			15853 => std_logic_vector(to_unsigned( 173,8)),
			15854 => std_logic_vector(to_unsigned( 75,8)),
			15855 => std_logic_vector(to_unsigned( 64,8)),
			15856 => std_logic_vector(to_unsigned( 43,8)),
			15857 => std_logic_vector(to_unsigned( 75,8)),
			15858 => std_logic_vector(to_unsigned( 214,8)),
			15859 => std_logic_vector(to_unsigned( 210,8)),
			15860 => std_logic_vector(to_unsigned( 104,8)),
			15861 => std_logic_vector(to_unsigned( 135,8)),
			15862 => std_logic_vector(to_unsigned( 199,8)),
			15863 => std_logic_vector(to_unsigned( 218,8)),
			15864 => std_logic_vector(to_unsigned( 81,8)),
			15865 => std_logic_vector(to_unsigned( 69,8)),
			15866 => std_logic_vector(to_unsigned( 94,8)),
			15867 => std_logic_vector(to_unsigned( 130,8)),
			15868 => std_logic_vector(to_unsigned( 50,8)),
			15869 => std_logic_vector(to_unsigned( 231,8)),
			15870 => std_logic_vector(to_unsigned( 126,8)),
			15871 => std_logic_vector(to_unsigned( 245,8)),
			15872 => std_logic_vector(to_unsigned( 229,8)),
			15873 => std_logic_vector(to_unsigned( 236,8)),
			15874 => std_logic_vector(to_unsigned( 175,8)),
			15875 => std_logic_vector(to_unsigned( 212,8)),
			15876 => std_logic_vector(to_unsigned( 64,8)),
			15877 => std_logic_vector(to_unsigned( 248,8)),
			15878 => std_logic_vector(to_unsigned( 17,8)),
			15879 => std_logic_vector(to_unsigned( 46,8)),
			15880 => std_logic_vector(to_unsigned( 245,8)),
			15881 => std_logic_vector(to_unsigned( 24,8)),
			15882 => std_logic_vector(to_unsigned( 236,8)),
			15883 => std_logic_vector(to_unsigned( 60,8)),
			15884 => std_logic_vector(to_unsigned( 237,8)),
			15885 => std_logic_vector(to_unsigned( 22,8)),
			15886 => std_logic_vector(to_unsigned( 249,8)),
			15887 => std_logic_vector(to_unsigned( 119,8)),
			15888 => std_logic_vector(to_unsigned( 122,8)),
			15889 => std_logic_vector(to_unsigned( 209,8)),
			15890 => std_logic_vector(to_unsigned( 18,8)),
			15891 => std_logic_vector(to_unsigned( 80,8)),
			15892 => std_logic_vector(to_unsigned( 51,8)),
			15893 => std_logic_vector(to_unsigned( 71,8)),
			15894 => std_logic_vector(to_unsigned( 232,8)),
			15895 => std_logic_vector(to_unsigned( 26,8)),
			15896 => std_logic_vector(to_unsigned( 157,8)),
			15897 => std_logic_vector(to_unsigned( 21,8)),
			15898 => std_logic_vector(to_unsigned( 236,8)),
			15899 => std_logic_vector(to_unsigned( 27,8)),
			15900 => std_logic_vector(to_unsigned( 47,8)),
			15901 => std_logic_vector(to_unsigned( 136,8)),
			15902 => std_logic_vector(to_unsigned( 122,8)),
			15903 => std_logic_vector(to_unsigned( 255,8)),
			15904 => std_logic_vector(to_unsigned( 244,8)),
			15905 => std_logic_vector(to_unsigned( 26,8)),
			15906 => std_logic_vector(to_unsigned( 164,8)),
			15907 => std_logic_vector(to_unsigned( 86,8)),
			15908 => std_logic_vector(to_unsigned( 199,8)),
			15909 => std_logic_vector(to_unsigned( 127,8)),
			15910 => std_logic_vector(to_unsigned( 28,8)),
			15911 => std_logic_vector(to_unsigned( 239,8)),
			15912 => std_logic_vector(to_unsigned( 112,8)),
			15913 => std_logic_vector(to_unsigned( 174,8)),
			15914 => std_logic_vector(to_unsigned( 178,8)),
			15915 => std_logic_vector(to_unsigned( 214,8)),
			15916 => std_logic_vector(to_unsigned( 143,8)),
			15917 => std_logic_vector(to_unsigned( 18,8)),
			15918 => std_logic_vector(to_unsigned( 44,8)),
			15919 => std_logic_vector(to_unsigned( 96,8)),
			15920 => std_logic_vector(to_unsigned( 12,8)),
			15921 => std_logic_vector(to_unsigned( 24,8)),
			15922 => std_logic_vector(to_unsigned( 85,8)),
			15923 => std_logic_vector(to_unsigned( 79,8)),
			15924 => std_logic_vector(to_unsigned( 99,8)),
			15925 => std_logic_vector(to_unsigned( 48,8)),
			15926 => std_logic_vector(to_unsigned( 163,8)),
			15927 => std_logic_vector(to_unsigned( 116,8)),
			15928 => std_logic_vector(to_unsigned( 108,8)),
			15929 => std_logic_vector(to_unsigned( 159,8)),
			15930 => std_logic_vector(to_unsigned( 105,8)),
			15931 => std_logic_vector(to_unsigned( 112,8)),
			15932 => std_logic_vector(to_unsigned( 152,8)),
			15933 => std_logic_vector(to_unsigned( 224,8)),
			15934 => std_logic_vector(to_unsigned( 234,8)),
			15935 => std_logic_vector(to_unsigned( 54,8)),
			15936 => std_logic_vector(to_unsigned( 74,8)),
			15937 => std_logic_vector(to_unsigned( 237,8)),
			15938 => std_logic_vector(to_unsigned( 84,8)),
			15939 => std_logic_vector(to_unsigned( 165,8)),
			15940 => std_logic_vector(to_unsigned( 168,8)),
			15941 => std_logic_vector(to_unsigned( 15,8)),
			15942 => std_logic_vector(to_unsigned( 180,8)),
			15943 => std_logic_vector(to_unsigned( 108,8)),
			15944 => std_logic_vector(to_unsigned( 68,8)),
			15945 => std_logic_vector(to_unsigned( 68,8)),
			15946 => std_logic_vector(to_unsigned( 71,8)),
			15947 => std_logic_vector(to_unsigned( 171,8)),
			15948 => std_logic_vector(to_unsigned( 106,8)),
			15949 => std_logic_vector(to_unsigned( 17,8)),
			15950 => std_logic_vector(to_unsigned( 201,8)),
			15951 => std_logic_vector(to_unsigned( 245,8)),
			15952 => std_logic_vector(to_unsigned( 116,8)),
			15953 => std_logic_vector(to_unsigned( 227,8)),
			15954 => std_logic_vector(to_unsigned( 232,8)),
			15955 => std_logic_vector(to_unsigned( 29,8)),
			15956 => std_logic_vector(to_unsigned( 191,8)),
			15957 => std_logic_vector(to_unsigned( 81,8)),
			15958 => std_logic_vector(to_unsigned( 59,8)),
			15959 => std_logic_vector(to_unsigned( 122,8)),
			15960 => std_logic_vector(to_unsigned( 205,8)),
			15961 => std_logic_vector(to_unsigned( 154,8)),
			15962 => std_logic_vector(to_unsigned( 7,8)),
			15963 => std_logic_vector(to_unsigned( 64,8)),
			15964 => std_logic_vector(to_unsigned( 47,8)),
			15965 => std_logic_vector(to_unsigned( 87,8)),
			15966 => std_logic_vector(to_unsigned( 201,8)),
			15967 => std_logic_vector(to_unsigned( 126,8)),
			15968 => std_logic_vector(to_unsigned( 114,8)),
			15969 => std_logic_vector(to_unsigned( 202,8)),
			15970 => std_logic_vector(to_unsigned( 213,8)),
			15971 => std_logic_vector(to_unsigned( 167,8)),
			15972 => std_logic_vector(to_unsigned( 75,8)),
			15973 => std_logic_vector(to_unsigned( 51,8)),
			15974 => std_logic_vector(to_unsigned( 206,8)),
			15975 => std_logic_vector(to_unsigned( 6,8)),
			15976 => std_logic_vector(to_unsigned( 129,8)),
			15977 => std_logic_vector(to_unsigned( 113,8)),
			15978 => std_logic_vector(to_unsigned( 127,8)),
			15979 => std_logic_vector(to_unsigned( 45,8)),
			15980 => std_logic_vector(to_unsigned( 231,8)),
			15981 => std_logic_vector(to_unsigned( 11,8)),
			15982 => std_logic_vector(to_unsigned( 33,8)),
			15983 => std_logic_vector(to_unsigned( 36,8)),
			15984 => std_logic_vector(to_unsigned( 128,8)),
			15985 => std_logic_vector(to_unsigned( 123,8)),
			15986 => std_logic_vector(to_unsigned( 142,8)),
			15987 => std_logic_vector(to_unsigned( 182,8)),
			15988 => std_logic_vector(to_unsigned( 168,8)),
			15989 => std_logic_vector(to_unsigned( 97,8)),
			15990 => std_logic_vector(to_unsigned( 156,8)),
			15991 => std_logic_vector(to_unsigned( 91,8)),
			15992 => std_logic_vector(to_unsigned( 156,8)),
			15993 => std_logic_vector(to_unsigned( 43,8)),
			15994 => std_logic_vector(to_unsigned( 238,8)),
			15995 => std_logic_vector(to_unsigned( 174,8)),
			15996 => std_logic_vector(to_unsigned( 156,8)),
			15997 => std_logic_vector(to_unsigned( 225,8)),
			15998 => std_logic_vector(to_unsigned( 119,8)),
			15999 => std_logic_vector(to_unsigned( 31,8)),
			16000 => std_logic_vector(to_unsigned( 187,8)),
			16001 => std_logic_vector(to_unsigned( 250,8)),
			16002 => std_logic_vector(to_unsigned( 135,8)),
			16003 => std_logic_vector(to_unsigned( 59,8)),
			16004 => std_logic_vector(to_unsigned( 90,8)),
			16005 => std_logic_vector(to_unsigned( 75,8)),
			16006 => std_logic_vector(to_unsigned( 219,8)),
			16007 => std_logic_vector(to_unsigned( 55,8)),
			16008 => std_logic_vector(to_unsigned( 91,8)),
			16009 => std_logic_vector(to_unsigned( 96,8)),
			16010 => std_logic_vector(to_unsigned( 178,8)),
			16011 => std_logic_vector(to_unsigned( 66,8)),
			16012 => std_logic_vector(to_unsigned( 107,8)),
			16013 => std_logic_vector(to_unsigned( 73,8)),
			16014 => std_logic_vector(to_unsigned( 52,8)),
			16015 => std_logic_vector(to_unsigned( 233,8)),
			16016 => std_logic_vector(to_unsigned( 146,8)),
			16017 => std_logic_vector(to_unsigned( 141,8)),
			16018 => std_logic_vector(to_unsigned( 136,8)),
			16019 => std_logic_vector(to_unsigned( 7,8)),
			16020 => std_logic_vector(to_unsigned( 10,8)),
			16021 => std_logic_vector(to_unsigned( 239,8)),
			16022 => std_logic_vector(to_unsigned( 213,8)),
			16023 => std_logic_vector(to_unsigned( 253,8)),
			16024 => std_logic_vector(to_unsigned( 7,8)),
			16025 => std_logic_vector(to_unsigned( 230,8)),
			16026 => std_logic_vector(to_unsigned( 33,8)),
			16027 => std_logic_vector(to_unsigned( 160,8)),
			16028 => std_logic_vector(to_unsigned( 145,8)),
			16029 => std_logic_vector(to_unsigned( 210,8)),
			16030 => std_logic_vector(to_unsigned( 20,8)),
			16031 => std_logic_vector(to_unsigned( 182,8)),
			16032 => std_logic_vector(to_unsigned( 33,8)),
			16033 => std_logic_vector(to_unsigned( 251,8)),
			16034 => std_logic_vector(to_unsigned( 1,8)),
			16035 => std_logic_vector(to_unsigned( 89,8)),
			16036 => std_logic_vector(to_unsigned( 34,8)),
			16037 => std_logic_vector(to_unsigned( 122,8)),
			16038 => std_logic_vector(to_unsigned( 111,8)),
			16039 => std_logic_vector(to_unsigned( 29,8)),
			16040 => std_logic_vector(to_unsigned( 148,8)),
			16041 => std_logic_vector(to_unsigned( 243,8)),
			16042 => std_logic_vector(to_unsigned( 246,8)),
			16043 => std_logic_vector(to_unsigned( 171,8)),
			16044 => std_logic_vector(to_unsigned( 183,8)),
			16045 => std_logic_vector(to_unsigned( 231,8)),
			16046 => std_logic_vector(to_unsigned( 137,8)),
			16047 => std_logic_vector(to_unsigned( 95,8)),
			16048 => std_logic_vector(to_unsigned( 181,8)),
			16049 => std_logic_vector(to_unsigned( 64,8)),
			16050 => std_logic_vector(to_unsigned( 113,8)),
			16051 => std_logic_vector(to_unsigned( 40,8)),
			16052 => std_logic_vector(to_unsigned( 212,8)),
			16053 => std_logic_vector(to_unsigned( 8,8)),
			16054 => std_logic_vector(to_unsigned( 76,8)),
			16055 => std_logic_vector(to_unsigned( 80,8)),
			16056 => std_logic_vector(to_unsigned( 40,8)),
			16057 => std_logic_vector(to_unsigned( 71,8)),
			16058 => std_logic_vector(to_unsigned( 89,8)),
			16059 => std_logic_vector(to_unsigned( 193,8)),
			16060 => std_logic_vector(to_unsigned( 227,8)),
			16061 => std_logic_vector(to_unsigned( 167,8)),
			16062 => std_logic_vector(to_unsigned( 242,8)),
			16063 => std_logic_vector(to_unsigned( 72,8)),
			16064 => std_logic_vector(to_unsigned( 225,8)),
			16065 => std_logic_vector(to_unsigned( 103,8)),
			16066 => std_logic_vector(to_unsigned( 250,8)),
			16067 => std_logic_vector(to_unsigned( 138,8)),
			16068 => std_logic_vector(to_unsigned( 173,8)),
			16069 => std_logic_vector(to_unsigned( 159,8)),
			16070 => std_logic_vector(to_unsigned( 53,8)),
			16071 => std_logic_vector(to_unsigned( 33,8)),
			16072 => std_logic_vector(to_unsigned( 237,8)),
			16073 => std_logic_vector(to_unsigned( 151,8)),
			16074 => std_logic_vector(to_unsigned( 50,8)),
			16075 => std_logic_vector(to_unsigned( 141,8)),
			16076 => std_logic_vector(to_unsigned( 130,8)),
			16077 => std_logic_vector(to_unsigned( 94,8)),
			16078 => std_logic_vector(to_unsigned( 68,8)),
			16079 => std_logic_vector(to_unsigned( 144,8)),
			16080 => std_logic_vector(to_unsigned( 30,8)),
			16081 => std_logic_vector(to_unsigned( 102,8)),
			16082 => std_logic_vector(to_unsigned( 236,8)),
			16083 => std_logic_vector(to_unsigned( 52,8)),
			16084 => std_logic_vector(to_unsigned( 191,8)),
			16085 => std_logic_vector(to_unsigned( 12,8)),
			16086 => std_logic_vector(to_unsigned( 74,8)),
			16087 => std_logic_vector(to_unsigned( 162,8)),
			16088 => std_logic_vector(to_unsigned( 127,8)),
			16089 => std_logic_vector(to_unsigned( 148,8)),
			16090 => std_logic_vector(to_unsigned( 232,8)),
			16091 => std_logic_vector(to_unsigned( 181,8)),
			16092 => std_logic_vector(to_unsigned( 196,8)),
			16093 => std_logic_vector(to_unsigned( 26,8)),
			16094 => std_logic_vector(to_unsigned( 22,8)),
			16095 => std_logic_vector(to_unsigned( 114,8)),
			16096 => std_logic_vector(to_unsigned( 210,8)),
			16097 => std_logic_vector(to_unsigned( 19,8)),
			16098 => std_logic_vector(to_unsigned( 37,8)),
			16099 => std_logic_vector(to_unsigned( 151,8)),
			16100 => std_logic_vector(to_unsigned( 148,8)),
			16101 => std_logic_vector(to_unsigned( 215,8)),
			16102 => std_logic_vector(to_unsigned( 209,8)),
			16103 => std_logic_vector(to_unsigned( 222,8)),
			16104 => std_logic_vector(to_unsigned( 188,8)),
			16105 => std_logic_vector(to_unsigned( 193,8)),
			16106 => std_logic_vector(to_unsigned( 152,8)),
			16107 => std_logic_vector(to_unsigned( 108,8)),
			16108 => std_logic_vector(to_unsigned( 157,8)),
			16109 => std_logic_vector(to_unsigned( 44,8)),
			16110 => std_logic_vector(to_unsigned( 180,8)),
			16111 => std_logic_vector(to_unsigned( 190,8)),
			16112 => std_logic_vector(to_unsigned( 129,8)),
			16113 => std_logic_vector(to_unsigned( 139,8)),
			16114 => std_logic_vector(to_unsigned( 178,8)),
			16115 => std_logic_vector(to_unsigned( 10,8)),
			16116 => std_logic_vector(to_unsigned( 231,8)),
			16117 => std_logic_vector(to_unsigned( 232,8)),
			16118 => std_logic_vector(to_unsigned( 38,8)),
			16119 => std_logic_vector(to_unsigned( 216,8)),
			16120 => std_logic_vector(to_unsigned( 59,8)),
			16121 => std_logic_vector(to_unsigned( 108,8)),
			16122 => std_logic_vector(to_unsigned( 241,8)),
			16123 => std_logic_vector(to_unsigned( 216,8)),
			16124 => std_logic_vector(to_unsigned( 96,8)),
			16125 => std_logic_vector(to_unsigned( 82,8)),
			16126 => std_logic_vector(to_unsigned( 225,8)),
			16127 => std_logic_vector(to_unsigned( 122,8)),
			16128 => std_logic_vector(to_unsigned( 60,8)),
			16129 => std_logic_vector(to_unsigned( 68,8)),
			16130 => std_logic_vector(to_unsigned( 207,8)),
			16131 => std_logic_vector(to_unsigned( 246,8)),
			16132 => std_logic_vector(to_unsigned( 111,8)),
			16133 => std_logic_vector(to_unsigned( 80,8)),
			16134 => std_logic_vector(to_unsigned( 252,8)),
			16135 => std_logic_vector(to_unsigned( 154,8)),
			16136 => std_logic_vector(to_unsigned( 194,8)),
			16137 => std_logic_vector(to_unsigned( 111,8)),
			16138 => std_logic_vector(to_unsigned( 29,8)),
			16139 => std_logic_vector(to_unsigned( 12,8)),
			16140 => std_logic_vector(to_unsigned( 68,8)),
			16141 => std_logic_vector(to_unsigned( 197,8)),
			16142 => std_logic_vector(to_unsigned( 34,8)),
			16143 => std_logic_vector(to_unsigned( 6,8)),
			16144 => std_logic_vector(to_unsigned( 154,8)),
			16145 => std_logic_vector(to_unsigned( 144,8)),
			16146 => std_logic_vector(to_unsigned( 181,8)),
			16147 => std_logic_vector(to_unsigned( 252,8)),
			16148 => std_logic_vector(to_unsigned( 66,8)),
			16149 => std_logic_vector(to_unsigned( 42,8)),
			16150 => std_logic_vector(to_unsigned( 20,8)),
			16151 => std_logic_vector(to_unsigned( 0,8)),
			16152 => std_logic_vector(to_unsigned( 39,8)),
			16153 => std_logic_vector(to_unsigned( 245,8)),
			16154 => std_logic_vector(to_unsigned( 250,8)),
			16155 => std_logic_vector(to_unsigned( 230,8)),
			16156 => std_logic_vector(to_unsigned( 22,8)),
			16157 => std_logic_vector(to_unsigned( 10,8)),
			16158 => std_logic_vector(to_unsigned( 52,8)),
			16159 => std_logic_vector(to_unsigned( 127,8)),
			16160 => std_logic_vector(to_unsigned( 189,8)),
			16161 => std_logic_vector(to_unsigned( 22,8)),
			16162 => std_logic_vector(to_unsigned( 247,8)),
			16163 => std_logic_vector(to_unsigned( 228,8)),
			16164 => std_logic_vector(to_unsigned( 64,8)),
			16165 => std_logic_vector(to_unsigned( 239,8)),
			16166 => std_logic_vector(to_unsigned( 183,8)),
			16167 => std_logic_vector(to_unsigned( 109,8)),
			16168 => std_logic_vector(to_unsigned( 97,8)),
			16169 => std_logic_vector(to_unsigned( 35,8)),
			16170 => std_logic_vector(to_unsigned( 220,8)),
			16171 => std_logic_vector(to_unsigned( 230,8)),
			16172 => std_logic_vector(to_unsigned( 172,8)),
			16173 => std_logic_vector(to_unsigned( 70,8)),
			16174 => std_logic_vector(to_unsigned( 32,8)),
			16175 => std_logic_vector(to_unsigned( 145,8)),
			16176 => std_logic_vector(to_unsigned( 87,8)),
			16177 => std_logic_vector(to_unsigned( 249,8)),
			16178 => std_logic_vector(to_unsigned( 22,8)),
			16179 => std_logic_vector(to_unsigned( 203,8)),
			16180 => std_logic_vector(to_unsigned( 234,8)),
			16181 => std_logic_vector(to_unsigned( 130,8)),
			16182 => std_logic_vector(to_unsigned( 210,8)),
			16183 => std_logic_vector(to_unsigned( 2,8)),
			16184 => std_logic_vector(to_unsigned( 159,8)),
			16185 => std_logic_vector(to_unsigned( 192,8)),
			16186 => std_logic_vector(to_unsigned( 105,8)),
			16187 => std_logic_vector(to_unsigned( 103,8)),
			16188 => std_logic_vector(to_unsigned( 74,8)),
			16189 => std_logic_vector(to_unsigned( 82,8)),
			16190 => std_logic_vector(to_unsigned( 160,8)),
			16191 => std_logic_vector(to_unsigned( 135,8)),
			16192 => std_logic_vector(to_unsigned( 140,8)),
			16193 => std_logic_vector(to_unsigned( 251,8)),
			16194 => std_logic_vector(to_unsigned( 202,8)),
			16195 => std_logic_vector(to_unsigned( 114,8)),
			16196 => std_logic_vector(to_unsigned( 213,8)),
			16197 => std_logic_vector(to_unsigned( 154,8)),
			16198 => std_logic_vector(to_unsigned( 79,8)),
			16199 => std_logic_vector(to_unsigned( 201,8)),
			16200 => std_logic_vector(to_unsigned( 229,8)),
			16201 => std_logic_vector(to_unsigned( 67,8)),
			16202 => std_logic_vector(to_unsigned( 69,8)),
			16203 => std_logic_vector(to_unsigned( 163,8)),
			16204 => std_logic_vector(to_unsigned( 17,8)),
			16205 => std_logic_vector(to_unsigned( 17,8)),
			16206 => std_logic_vector(to_unsigned( 213,8)),
			16207 => std_logic_vector(to_unsigned( 225,8)),
			16208 => std_logic_vector(to_unsigned( 96,8)),
			16209 => std_logic_vector(to_unsigned( 24,8)),
			16210 => std_logic_vector(to_unsigned( 43,8)),
			16211 => std_logic_vector(to_unsigned( 205,8)),
			16212 => std_logic_vector(to_unsigned( 85,8)),
			16213 => std_logic_vector(to_unsigned( 16,8)),
			16214 => std_logic_vector(to_unsigned( 182,8)),
			16215 => std_logic_vector(to_unsigned( 227,8)),
			16216 => std_logic_vector(to_unsigned( 217,8)),
			16217 => std_logic_vector(to_unsigned( 133,8)),
			16218 => std_logic_vector(to_unsigned( 241,8)),
			16219 => std_logic_vector(to_unsigned( 128,8)),
			16220 => std_logic_vector(to_unsigned( 196,8)),
			16221 => std_logic_vector(to_unsigned( 27,8)),
			16222 => std_logic_vector(to_unsigned( 28,8)),
			16223 => std_logic_vector(to_unsigned( 139,8)),
			16224 => std_logic_vector(to_unsigned( 168,8)),
			16225 => std_logic_vector(to_unsigned( 242,8)),
			16226 => std_logic_vector(to_unsigned( 202,8)),
			16227 => std_logic_vector(to_unsigned( 228,8)),
			16228 => std_logic_vector(to_unsigned( 90,8)),
			16229 => std_logic_vector(to_unsigned( 148,8)),
			16230 => std_logic_vector(to_unsigned( 71,8)),
			16231 => std_logic_vector(to_unsigned( 22,8)),
			16232 => std_logic_vector(to_unsigned( 32,8)),
			16233 => std_logic_vector(to_unsigned( 230,8)),
			16234 => std_logic_vector(to_unsigned( 20,8)),
			16235 => std_logic_vector(to_unsigned( 96,8)),
			16236 => std_logic_vector(to_unsigned( 230,8)),
			16237 => std_logic_vector(to_unsigned( 10,8)),
			16238 => std_logic_vector(to_unsigned( 0,8)),
			16239 => std_logic_vector(to_unsigned( 120,8)),
			16240 => std_logic_vector(to_unsigned( 157,8)),
			16241 => std_logic_vector(to_unsigned( 92,8)),
			16242 => std_logic_vector(to_unsigned( 169,8)),
			16243 => std_logic_vector(to_unsigned( 172,8)),
			16244 => std_logic_vector(to_unsigned( 83,8)),
			16245 => std_logic_vector(to_unsigned( 252,8)),
			16246 => std_logic_vector(to_unsigned( 6,8)),
			16247 => std_logic_vector(to_unsigned( 100,8)),
			16248 => std_logic_vector(to_unsigned( 96,8)),
			16249 => std_logic_vector(to_unsigned( 224,8)),
			16250 => std_logic_vector(to_unsigned( 18,8)),
			16251 => std_logic_vector(to_unsigned( 202,8)),
			16252 => std_logic_vector(to_unsigned( 147,8)),
			16253 => std_logic_vector(to_unsigned( 121,8)),
			16254 => std_logic_vector(to_unsigned( 165,8)),
			16255 => std_logic_vector(to_unsigned( 61,8)),
			16256 => std_logic_vector(to_unsigned( 76,8)),
			16257 => std_logic_vector(to_unsigned( 83,8)),
			16258 => std_logic_vector(to_unsigned( 178,8)),
			16259 => std_logic_vector(to_unsigned( 145,8)),
			16260 => std_logic_vector(to_unsigned( 59,8)),
			16261 => std_logic_vector(to_unsigned( 33,8)),
			16262 => std_logic_vector(to_unsigned( 29,8)),
			16263 => std_logic_vector(to_unsigned( 208,8)),
			16264 => std_logic_vector(to_unsigned( 9,8)),
			16265 => std_logic_vector(to_unsigned( 225,8)),
			16266 => std_logic_vector(to_unsigned( 94,8)),
			16267 => std_logic_vector(to_unsigned( 212,8)),
			16268 => std_logic_vector(to_unsigned( 195,8)),
			16269 => std_logic_vector(to_unsigned( 48,8)),
			16270 => std_logic_vector(to_unsigned( 197,8)),
			16271 => std_logic_vector(to_unsigned( 73,8)),
			16272 => std_logic_vector(to_unsigned( 190,8)),
			16273 => std_logic_vector(to_unsigned( 4,8)),
			16274 => std_logic_vector(to_unsigned( 93,8)),
			16275 => std_logic_vector(to_unsigned( 86,8)),
			16276 => std_logic_vector(to_unsigned( 89,8)),
			16277 => std_logic_vector(to_unsigned( 38,8)),
			16278 => std_logic_vector(to_unsigned( 199,8)),
			16279 => std_logic_vector(to_unsigned( 26,8)),
			16280 => std_logic_vector(to_unsigned( 181,8)),
			16281 => std_logic_vector(to_unsigned( 135,8)),
			16282 => std_logic_vector(to_unsigned( 225,8)),
			16283 => std_logic_vector(to_unsigned( 37,8)),
			16284 => std_logic_vector(to_unsigned( 93,8)),
			16285 => std_logic_vector(to_unsigned( 226,8)),
			16286 => std_logic_vector(to_unsigned( 121,8)),
			16287 => std_logic_vector(to_unsigned( 253,8)),
			16288 => std_logic_vector(to_unsigned( 132,8)),
			16289 => std_logic_vector(to_unsigned( 185,8)),
			16290 => std_logic_vector(to_unsigned( 150,8)),
			16291 => std_logic_vector(to_unsigned( 161,8)),
			16292 => std_logic_vector(to_unsigned( 227,8)),
			16293 => std_logic_vector(to_unsigned( 202,8)),
			16294 => std_logic_vector(to_unsigned( 78,8)),
			16295 => std_logic_vector(to_unsigned( 69,8)),
			16296 => std_logic_vector(to_unsigned( 208,8)),
			16297 => std_logic_vector(to_unsigned( 33,8)),
			16298 => std_logic_vector(to_unsigned( 188,8)),
			16299 => std_logic_vector(to_unsigned( 41,8)),
			16300 => std_logic_vector(to_unsigned( 57,8)),
			16301 => std_logic_vector(to_unsigned( 250,8)),
			16302 => std_logic_vector(to_unsigned( 210,8)),
			16303 => std_logic_vector(to_unsigned( 37,8)),
			16304 => std_logic_vector(to_unsigned( 117,8)),
			16305 => std_logic_vector(to_unsigned( 35,8)),
			16306 => std_logic_vector(to_unsigned( 60,8)),
			16307 => std_logic_vector(to_unsigned( 80,8)),
			16308 => std_logic_vector(to_unsigned( 255,8)),
			16309 => std_logic_vector(to_unsigned( 50,8)),
			16310 => std_logic_vector(to_unsigned( 192,8)),
			16311 => std_logic_vector(to_unsigned( 89,8)),
			16312 => std_logic_vector(to_unsigned( 245,8)),
			16313 => std_logic_vector(to_unsigned( 93,8)),
			16314 => std_logic_vector(to_unsigned( 197,8)),
			16315 => std_logic_vector(to_unsigned( 130,8)),
			16316 => std_logic_vector(to_unsigned( 18,8)),
			16317 => std_logic_vector(to_unsigned( 4,8)),
			16318 => std_logic_vector(to_unsigned( 197,8)),
			16319 => std_logic_vector(to_unsigned( 217,8)),
			16320 => std_logic_vector(to_unsigned( 225,8)),
			16321 => std_logic_vector(to_unsigned( 157,8)),
			16322 => std_logic_vector(to_unsigned( 149,8)),
			16323 => std_logic_vector(to_unsigned( 11,8)),
			16324 => std_logic_vector(to_unsigned( 46,8)),
			16325 => std_logic_vector(to_unsigned( 163,8)),
			16326 => std_logic_vector(to_unsigned( 67,8)),
			16327 => std_logic_vector(to_unsigned( 21,8)),
			16328 => std_logic_vector(to_unsigned( 208,8)),
			16329 => std_logic_vector(to_unsigned( 171,8)),
			16330 => std_logic_vector(to_unsigned( 178,8)),
			16331 => std_logic_vector(to_unsigned( 221,8)),
			16332 => std_logic_vector(to_unsigned( 223,8)),
			16333 => std_logic_vector(to_unsigned( 160,8)),
			16334 => std_logic_vector(to_unsigned( 149,8)),
			16335 => std_logic_vector(to_unsigned( 47,8)),
			16336 => std_logic_vector(to_unsigned( 164,8)),
			16337 => std_logic_vector(to_unsigned( 180,8)),
			16338 => std_logic_vector(to_unsigned( 185,8)),
			16339 => std_logic_vector(to_unsigned( 166,8)),
			16340 => std_logic_vector(to_unsigned( 211,8)),
			16341 => std_logic_vector(to_unsigned( 41,8)),
			16342 => std_logic_vector(to_unsigned( 140,8)),
			16343 => std_logic_vector(to_unsigned( 10,8)),
			16344 => std_logic_vector(to_unsigned( 181,8)),
			16345 => std_logic_vector(to_unsigned( 7,8)),
			16346 => std_logic_vector(to_unsigned( 54,8)),
			16347 => std_logic_vector(to_unsigned( 30,8)),
			16348 => std_logic_vector(to_unsigned( 30,8)),
			16349 => std_logic_vector(to_unsigned( 179,8)),
			16350 => std_logic_vector(to_unsigned( 30,8)),
			16351 => std_logic_vector(to_unsigned( 212,8)),
			16352 => std_logic_vector(to_unsigned( 149,8)),
			16353 => std_logic_vector(to_unsigned( 101,8)),
			16354 => std_logic_vector(to_unsigned( 49,8)),
			16355 => std_logic_vector(to_unsigned( 33,8)),
			16356 => std_logic_vector(to_unsigned( 186,8)),
			16357 => std_logic_vector(to_unsigned( 68,8)),
			16358 => std_logic_vector(to_unsigned( 79,8)),
			16359 => std_logic_vector(to_unsigned( 186,8)),
			16360 => std_logic_vector(to_unsigned( 101,8)),
			16361 => std_logic_vector(to_unsigned( 239,8)),
			16362 => std_logic_vector(to_unsigned( 63,8)),
			16363 => std_logic_vector(to_unsigned( 246,8)),
			16364 => std_logic_vector(to_unsigned( 46,8)),
			16365 => std_logic_vector(to_unsigned( 129,8)),
			16366 => std_logic_vector(to_unsigned( 212,8)),
			16367 => std_logic_vector(to_unsigned( 236,8)),
			16368 => std_logic_vector(to_unsigned( 208,8)),
			16369 => std_logic_vector(to_unsigned( 122,8)),
			16370 => std_logic_vector(to_unsigned( 191,8)),
			16371 => std_logic_vector(to_unsigned( 248,8)),
			16372 => std_logic_vector(to_unsigned( 234,8)),
			16373 => std_logic_vector(to_unsigned( 113,8)),
			16374 => std_logic_vector(to_unsigned( 122,8)),
			16375 => std_logic_vector(to_unsigned( 203,8)),
			16376 => std_logic_vector(to_unsigned( 233,8)),
			16377 => std_logic_vector(to_unsigned( 53,8)),
			16378 => std_logic_vector(to_unsigned( 196,8)),
			16379 => std_logic_vector(to_unsigned( 2,8)),
			16380 => std_logic_vector(to_unsigned( 162,8)),
			16381 => std_logic_vector(to_unsigned( 167,8)),
			16382 => std_logic_vector(to_unsigned( 229,8)),
			16383 => std_logic_vector(to_unsigned( 29,8)),
			16384 => std_logic_vector(to_unsigned( 235,8)),
			16385 => std_logic_vector(to_unsigned( 105,8)),
			others => (others => '0'));


			 -- Expected Output  6 -> 0                         
			 -- Expected Output  7 -> 255                         
			 -- Expected Output  8 -> 64                         
			 -- Expected Output  9 -> 172                         

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;


test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;

    -- Immagine originale =  [46, 131, 62, 89]  
    -- Immagine di output =  [0, 255, 64, 172]  
    
	assert RAM(16386) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16386))))  severity failure;
	assert RAM(16387) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16387))))  severity failure;
	assert RAM(16388) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16388))))  severity failure;
	assert RAM(16389) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16389))))  severity failure;
	assert RAM(16390) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16390))))  severity failure;
	assert RAM(16391) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16391))))  severity failure;
	assert RAM(16392) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16392))))  severity failure;
	assert RAM(16393) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16393))))  severity failure;
	assert RAM(16394) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16394))))  severity failure;
	assert RAM(16395) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16395))))  severity failure;
	assert RAM(16396) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16396))))  severity failure;
	assert RAM(16397) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16397))))  severity failure;
	assert RAM(16398) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16398))))  severity failure;
	assert RAM(16399) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16399))))  severity failure;
	assert RAM(16400) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16400))))  severity failure;
	assert RAM(16401) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16401))))  severity failure;
	assert RAM(16402) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(16402))))  severity failure;
	assert RAM(16403) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(16403))))  severity failure;
	assert RAM(16404) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16404))))  severity failure;
	assert RAM(16405) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(16405))))  severity failure;
	assert RAM(16406) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16406))))  severity failure;
	assert RAM(16407) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(16407))))  severity failure;
	assert RAM(16408) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(16408))))  severity failure;
	assert RAM(16409) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16409))))  severity failure;
	assert RAM(16410) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16410))))  severity failure;
	assert RAM(16411) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(16411))))  severity failure;
	assert RAM(16412) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16412))))  severity failure;
	assert RAM(16413) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16413))))  severity failure;
	assert RAM(16414) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(16414))))  severity failure;
	assert RAM(16415) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16415))))  severity failure;
	assert RAM(16416) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16416))))  severity failure;
	assert RAM(16417) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16417))))  severity failure;
	assert RAM(16418) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16418))))  severity failure;
	assert RAM(16419) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(16419))))  severity failure;
	assert RAM(16420) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16420))))  severity failure;
	assert RAM(16421) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(16421))))  severity failure;
	assert RAM(16422) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16422))))  severity failure;
	assert RAM(16423) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16423))))  severity failure;
	assert RAM(16424) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(16424))))  severity failure;
	assert RAM(16425) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16425))))  severity failure;
	assert RAM(16426) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16426))))  severity failure;
	assert RAM(16427) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(16427))))  severity failure;
	assert RAM(16428) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16428))))  severity failure;
	assert RAM(16429) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16429))))  severity failure;
	assert RAM(16430) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16430))))  severity failure;
	assert RAM(16431) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16431))))  severity failure;
	assert RAM(16432) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16432))))  severity failure;
	assert RAM(16433) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16433))))  severity failure;
	assert RAM(16434) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16434))))  severity failure;
	assert RAM(16435) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(16435))))  severity failure;
	assert RAM(16436) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(16436))))  severity failure;
	assert RAM(16437) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(16437))))  severity failure;
	assert RAM(16438) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(16438))))  severity failure;
	assert RAM(16439) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(16439))))  severity failure;
	assert RAM(16440) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16440))))  severity failure;
	assert RAM(16441) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16441))))  severity failure;
	assert RAM(16442) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16442))))  severity failure;
	assert RAM(16443) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16443))))  severity failure;
	assert RAM(16444) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16444))))  severity failure;
	assert RAM(16445) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16445))))  severity failure;
	assert RAM(16446) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16446))))  severity failure;
	assert RAM(16447) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16447))))  severity failure;
	assert RAM(16448) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(16448))))  severity failure;
	assert RAM(16449) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16449))))  severity failure;
	assert RAM(16450) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16450))))  severity failure;
	assert RAM(16451) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(16451))))  severity failure;
	assert RAM(16452) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16452))))  severity failure;
	assert RAM(16453) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16453))))  severity failure;
	assert RAM(16454) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(16454))))  severity failure;
	assert RAM(16455) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16455))))  severity failure;
	assert RAM(16456) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16456))))  severity failure;
	assert RAM(16457) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(16457))))  severity failure;
	assert RAM(16458) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16458))))  severity failure;
	assert RAM(16459) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(16459))))  severity failure;
	assert RAM(16460) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16460))))  severity failure;
	assert RAM(16461) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16461))))  severity failure;
	assert RAM(16462) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16462))))  severity failure;
	assert RAM(16463) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16463))))  severity failure;
	assert RAM(16464) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16464))))  severity failure;
	assert RAM(16465) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16465))))  severity failure;
	assert RAM(16466) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(16466))))  severity failure;
	assert RAM(16467) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16467))))  severity failure;
	assert RAM(16468) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16468))))  severity failure;
	assert RAM(16469) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16469))))  severity failure;
	assert RAM(16470) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16470))))  severity failure;
	assert RAM(16471) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(16471))))  severity failure;
	assert RAM(16472) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16472))))  severity failure;
	assert RAM(16473) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(16473))))  severity failure;
	assert RAM(16474) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(16474))))  severity failure;
	assert RAM(16475) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16475))))  severity failure;
	assert RAM(16476) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16476))))  severity failure;
	assert RAM(16477) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(16477))))  severity failure;
	assert RAM(16478) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16478))))  severity failure;
	assert RAM(16479) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16479))))  severity failure;
	assert RAM(16480) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16480))))  severity failure;
	assert RAM(16481) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16481))))  severity failure;
	assert RAM(16482) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16482))))  severity failure;
	assert RAM(16483) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16483))))  severity failure;
	assert RAM(16484) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16484))))  severity failure;
	assert RAM(16485) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(16485))))  severity failure;
	assert RAM(16486) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16486))))  severity failure;
	assert RAM(16487) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16487))))  severity failure;
	assert RAM(16488) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16488))))  severity failure;
	assert RAM(16489) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16489))))  severity failure;
	assert RAM(16490) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16490))))  severity failure;
	assert RAM(16491) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16491))))  severity failure;
	assert RAM(16492) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16492))))  severity failure;
	assert RAM(16493) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(16493))))  severity failure;
	assert RAM(16494) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(16494))))  severity failure;
	assert RAM(16495) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16495))))  severity failure;
	assert RAM(16496) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16496))))  severity failure;
	assert RAM(16497) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16497))))  severity failure;
	assert RAM(16498) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16498))))  severity failure;
	assert RAM(16499) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16499))))  severity failure;
	assert RAM(16500) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16500))))  severity failure;
	assert RAM(16501) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16501))))  severity failure;
	assert RAM(16502) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(16502))))  severity failure;
	assert RAM(16503) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16503))))  severity failure;
	assert RAM(16504) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16504))))  severity failure;
	assert RAM(16505) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16505))))  severity failure;
	assert RAM(16506) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16506))))  severity failure;
	assert RAM(16507) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16507))))  severity failure;
	assert RAM(16508) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(16508))))  severity failure;
	assert RAM(16509) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(16509))))  severity failure;
	assert RAM(16510) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16510))))  severity failure;
	assert RAM(16511) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16511))))  severity failure;
	assert RAM(16512) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(16512))))  severity failure;
	assert RAM(16513) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16513))))  severity failure;
	assert RAM(16514) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16514))))  severity failure;
	assert RAM(16515) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16515))))  severity failure;
	assert RAM(16516) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(16516))))  severity failure;
	assert RAM(16517) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16517))))  severity failure;
	assert RAM(16518) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(16518))))  severity failure;
	assert RAM(16519) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16519))))  severity failure;
	assert RAM(16520) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16520))))  severity failure;
	assert RAM(16521) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16521))))  severity failure;
	assert RAM(16522) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(16522))))  severity failure;
	assert RAM(16523) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16523))))  severity failure;
	assert RAM(16524) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(16524))))  severity failure;
	assert RAM(16525) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16525))))  severity failure;
	assert RAM(16526) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(16526))))  severity failure;
	assert RAM(16527) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(16527))))  severity failure;
	assert RAM(16528) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(16528))))  severity failure;
	assert RAM(16529) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16529))))  severity failure;
	assert RAM(16530) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(16530))))  severity failure;
	assert RAM(16531) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(16531))))  severity failure;
	assert RAM(16532) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16532))))  severity failure;
	assert RAM(16533) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16533))))  severity failure;
	assert RAM(16534) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(16534))))  severity failure;
	assert RAM(16535) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16535))))  severity failure;
	assert RAM(16536) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16536))))  severity failure;
	assert RAM(16537) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16537))))  severity failure;
	assert RAM(16538) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(16538))))  severity failure;
	assert RAM(16539) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16539))))  severity failure;
	assert RAM(16540) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16540))))  severity failure;
	assert RAM(16541) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16541))))  severity failure;
	assert RAM(16542) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16542))))  severity failure;
	assert RAM(16543) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16543))))  severity failure;
	assert RAM(16544) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(16544))))  severity failure;
	assert RAM(16545) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16545))))  severity failure;
	assert RAM(16546) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16546))))  severity failure;
	assert RAM(16547) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(16547))))  severity failure;
	assert RAM(16548) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16548))))  severity failure;
	assert RAM(16549) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16549))))  severity failure;
	assert RAM(16550) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(16550))))  severity failure;
	assert RAM(16551) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16551))))  severity failure;
	assert RAM(16552) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(16552))))  severity failure;
	assert RAM(16553) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(16553))))  severity failure;
	assert RAM(16554) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(16554))))  severity failure;
	assert RAM(16555) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16555))))  severity failure;
	assert RAM(16556) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16556))))  severity failure;
	assert RAM(16557) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16557))))  severity failure;
	assert RAM(16558) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16558))))  severity failure;
	assert RAM(16559) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16559))))  severity failure;
	assert RAM(16560) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(16560))))  severity failure;
	assert RAM(16561) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(16561))))  severity failure;
	assert RAM(16562) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16562))))  severity failure;
	assert RAM(16563) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16563))))  severity failure;
	assert RAM(16564) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(16564))))  severity failure;
	assert RAM(16565) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16565))))  severity failure;
	assert RAM(16566) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16566))))  severity failure;
	assert RAM(16567) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16567))))  severity failure;
	assert RAM(16568) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16568))))  severity failure;
	assert RAM(16569) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16569))))  severity failure;
	assert RAM(16570) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16570))))  severity failure;
	assert RAM(16571) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16571))))  severity failure;
	assert RAM(16572) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16572))))  severity failure;
	assert RAM(16573) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(16573))))  severity failure;
	assert RAM(16574) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16574))))  severity failure;
	assert RAM(16575) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16575))))  severity failure;
	assert RAM(16576) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16576))))  severity failure;
	assert RAM(16577) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16577))))  severity failure;
	assert RAM(16578) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16578))))  severity failure;
	assert RAM(16579) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16579))))  severity failure;
	assert RAM(16580) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16580))))  severity failure;
	assert RAM(16581) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(16581))))  severity failure;
	assert RAM(16582) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16582))))  severity failure;
	assert RAM(16583) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16583))))  severity failure;
	assert RAM(16584) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16584))))  severity failure;
	assert RAM(16585) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16585))))  severity failure;
	assert RAM(16586) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16586))))  severity failure;
	assert RAM(16587) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(16587))))  severity failure;
	assert RAM(16588) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16588))))  severity failure;
	assert RAM(16589) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16589))))  severity failure;
	assert RAM(16590) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(16590))))  severity failure;
	assert RAM(16591) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(16591))))  severity failure;
	assert RAM(16592) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16592))))  severity failure;
	assert RAM(16593) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16593))))  severity failure;
	assert RAM(16594) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16594))))  severity failure;
	assert RAM(16595) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(16595))))  severity failure;
	assert RAM(16596) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(16596))))  severity failure;
	assert RAM(16597) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16597))))  severity failure;
	assert RAM(16598) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16598))))  severity failure;
	assert RAM(16599) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(16599))))  severity failure;
	assert RAM(16600) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16600))))  severity failure;
	assert RAM(16601) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(16601))))  severity failure;
	assert RAM(16602) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16602))))  severity failure;
	assert RAM(16603) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16603))))  severity failure;
	assert RAM(16604) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16604))))  severity failure;
	assert RAM(16605) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(16605))))  severity failure;
	assert RAM(16606) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16606))))  severity failure;
	assert RAM(16607) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16607))))  severity failure;
	assert RAM(16608) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16608))))  severity failure;
	assert RAM(16609) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16609))))  severity failure;
	assert RAM(16610) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16610))))  severity failure;
	assert RAM(16611) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16611))))  severity failure;
	assert RAM(16612) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16612))))  severity failure;
	assert RAM(16613) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16613))))  severity failure;
	assert RAM(16614) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16614))))  severity failure;
	assert RAM(16615) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16615))))  severity failure;
	assert RAM(16616) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16616))))  severity failure;
	assert RAM(16617) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16617))))  severity failure;
	assert RAM(16618) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16618))))  severity failure;
	assert RAM(16619) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16619))))  severity failure;
	assert RAM(16620) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16620))))  severity failure;
	assert RAM(16621) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(16621))))  severity failure;
	assert RAM(16622) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16622))))  severity failure;
	assert RAM(16623) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(16623))))  severity failure;
	assert RAM(16624) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(16624))))  severity failure;
	assert RAM(16625) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16625))))  severity failure;
	assert RAM(16626) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(16626))))  severity failure;
	assert RAM(16627) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16627))))  severity failure;
	assert RAM(16628) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16628))))  severity failure;
	assert RAM(16629) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(16629))))  severity failure;
	assert RAM(16630) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(16630))))  severity failure;
	assert RAM(16631) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16631))))  severity failure;
	assert RAM(16632) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16632))))  severity failure;
	assert RAM(16633) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16633))))  severity failure;
	assert RAM(16634) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16634))))  severity failure;
	assert RAM(16635) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(16635))))  severity failure;
	assert RAM(16636) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16636))))  severity failure;
	assert RAM(16637) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(16637))))  severity failure;
	assert RAM(16638) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(16638))))  severity failure;
	assert RAM(16639) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16639))))  severity failure;
	assert RAM(16640) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(16640))))  severity failure;
	assert RAM(16641) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16641))))  severity failure;
	assert RAM(16642) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16642))))  severity failure;
	assert RAM(16643) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16643))))  severity failure;
	assert RAM(16644) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16644))))  severity failure;
	assert RAM(16645) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16645))))  severity failure;
	assert RAM(16646) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16646))))  severity failure;
	assert RAM(16647) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16647))))  severity failure;
	assert RAM(16648) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(16648))))  severity failure;
	assert RAM(16649) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16649))))  severity failure;
	assert RAM(16650) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16650))))  severity failure;
	assert RAM(16651) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16651))))  severity failure;
	assert RAM(16652) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16652))))  severity failure;
	assert RAM(16653) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16653))))  severity failure;
	assert RAM(16654) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16654))))  severity failure;
	assert RAM(16655) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16655))))  severity failure;
	assert RAM(16656) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16656))))  severity failure;
	assert RAM(16657) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(16657))))  severity failure;
	assert RAM(16658) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16658))))  severity failure;
	assert RAM(16659) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(16659))))  severity failure;
	assert RAM(16660) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(16660))))  severity failure;
	assert RAM(16661) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(16661))))  severity failure;
	assert RAM(16662) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16662))))  severity failure;
	assert RAM(16663) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16663))))  severity failure;
	assert RAM(16664) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16664))))  severity failure;
	assert RAM(16665) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16665))))  severity failure;
	assert RAM(16666) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(16666))))  severity failure;
	assert RAM(16667) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16667))))  severity failure;
	assert RAM(16668) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16668))))  severity failure;
	assert RAM(16669) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16669))))  severity failure;
	assert RAM(16670) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(16670))))  severity failure;
	assert RAM(16671) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16671))))  severity failure;
	assert RAM(16672) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(16672))))  severity failure;
	assert RAM(16673) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16673))))  severity failure;
	assert RAM(16674) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(16674))))  severity failure;
	assert RAM(16675) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16675))))  severity failure;
	assert RAM(16676) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(16676))))  severity failure;
	assert RAM(16677) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16677))))  severity failure;
	assert RAM(16678) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16678))))  severity failure;
	assert RAM(16679) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16679))))  severity failure;
	assert RAM(16680) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(16680))))  severity failure;
	assert RAM(16681) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16681))))  severity failure;
	assert RAM(16682) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16682))))  severity failure;
	assert RAM(16683) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(16683))))  severity failure;
	assert RAM(16684) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16684))))  severity failure;
	assert RAM(16685) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(16685))))  severity failure;
	assert RAM(16686) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(16686))))  severity failure;
	assert RAM(16687) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16687))))  severity failure;
	assert RAM(16688) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16688))))  severity failure;
	assert RAM(16689) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16689))))  severity failure;
	assert RAM(16690) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(16690))))  severity failure;
	assert RAM(16691) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16691))))  severity failure;
	assert RAM(16692) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16692))))  severity failure;
	assert RAM(16693) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(16693))))  severity failure;
	assert RAM(16694) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(16694))))  severity failure;
	assert RAM(16695) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(16695))))  severity failure;
	assert RAM(16696) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(16696))))  severity failure;
	assert RAM(16697) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(16697))))  severity failure;
	assert RAM(16698) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16698))))  severity failure;
	assert RAM(16699) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(16699))))  severity failure;
	assert RAM(16700) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16700))))  severity failure;
	assert RAM(16701) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16701))))  severity failure;
	assert RAM(16702) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16702))))  severity failure;
	assert RAM(16703) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16703))))  severity failure;
	assert RAM(16704) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16704))))  severity failure;
	assert RAM(16705) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(16705))))  severity failure;
	assert RAM(16706) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16706))))  severity failure;
	assert RAM(16707) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16707))))  severity failure;
	assert RAM(16708) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16708))))  severity failure;
	assert RAM(16709) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16709))))  severity failure;
	assert RAM(16710) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16710))))  severity failure;
	assert RAM(16711) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(16711))))  severity failure;
	assert RAM(16712) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16712))))  severity failure;
	assert RAM(16713) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(16713))))  severity failure;
	assert RAM(16714) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16714))))  severity failure;
	assert RAM(16715) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16715))))  severity failure;
	assert RAM(16716) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16716))))  severity failure;
	assert RAM(16717) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16717))))  severity failure;
	assert RAM(16718) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16718))))  severity failure;
	assert RAM(16719) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16719))))  severity failure;
	assert RAM(16720) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16720))))  severity failure;
	assert RAM(16721) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16721))))  severity failure;
	assert RAM(16722) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16722))))  severity failure;
	assert RAM(16723) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(16723))))  severity failure;
	assert RAM(16724) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16724))))  severity failure;
	assert RAM(16725) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16725))))  severity failure;
	assert RAM(16726) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16726))))  severity failure;
	assert RAM(16727) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16727))))  severity failure;
	assert RAM(16728) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(16728))))  severity failure;
	assert RAM(16729) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16729))))  severity failure;
	assert RAM(16730) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16730))))  severity failure;
	assert RAM(16731) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16731))))  severity failure;
	assert RAM(16732) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(16732))))  severity failure;
	assert RAM(16733) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(16733))))  severity failure;
	assert RAM(16734) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16734))))  severity failure;
	assert RAM(16735) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16735))))  severity failure;
	assert RAM(16736) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16736))))  severity failure;
	assert RAM(16737) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16737))))  severity failure;
	assert RAM(16738) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16738))))  severity failure;
	assert RAM(16739) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16739))))  severity failure;
	assert RAM(16740) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16740))))  severity failure;
	assert RAM(16741) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(16741))))  severity failure;
	assert RAM(16742) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16742))))  severity failure;
	assert RAM(16743) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16743))))  severity failure;
	assert RAM(16744) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16744))))  severity failure;
	assert RAM(16745) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16745))))  severity failure;
	assert RAM(16746) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(16746))))  severity failure;
	assert RAM(16747) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16747))))  severity failure;
	assert RAM(16748) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16748))))  severity failure;
	assert RAM(16749) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16749))))  severity failure;
	assert RAM(16750) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16750))))  severity failure;
	assert RAM(16751) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16751))))  severity failure;
	assert RAM(16752) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(16752))))  severity failure;
	assert RAM(16753) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16753))))  severity failure;
	assert RAM(16754) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(16754))))  severity failure;
	assert RAM(16755) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16755))))  severity failure;
	assert RAM(16756) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16756))))  severity failure;
	assert RAM(16757) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(16757))))  severity failure;
	assert RAM(16758) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16758))))  severity failure;
	assert RAM(16759) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16759))))  severity failure;
	assert RAM(16760) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16760))))  severity failure;
	assert RAM(16761) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16761))))  severity failure;
	assert RAM(16762) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16762))))  severity failure;
	assert RAM(16763) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16763))))  severity failure;
	assert RAM(16764) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16764))))  severity failure;
	assert RAM(16765) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16765))))  severity failure;
	assert RAM(16766) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16766))))  severity failure;
	assert RAM(16767) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16767))))  severity failure;
	assert RAM(16768) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16768))))  severity failure;
	assert RAM(16769) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(16769))))  severity failure;
	assert RAM(16770) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16770))))  severity failure;
	assert RAM(16771) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16771))))  severity failure;
	assert RAM(16772) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16772))))  severity failure;
	assert RAM(16773) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(16773))))  severity failure;
	assert RAM(16774) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(16774))))  severity failure;
	assert RAM(16775) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16775))))  severity failure;
	assert RAM(16776) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(16776))))  severity failure;
	assert RAM(16777) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16777))))  severity failure;
	assert RAM(16778) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16778))))  severity failure;
	assert RAM(16779) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16779))))  severity failure;
	assert RAM(16780) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(16780))))  severity failure;
	assert RAM(16781) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16781))))  severity failure;
	assert RAM(16782) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16782))))  severity failure;
	assert RAM(16783) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16783))))  severity failure;
	assert RAM(16784) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(16784))))  severity failure;
	assert RAM(16785) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(16785))))  severity failure;
	assert RAM(16786) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(16786))))  severity failure;
	assert RAM(16787) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16787))))  severity failure;
	assert RAM(16788) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16788))))  severity failure;
	assert RAM(16789) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16789))))  severity failure;
	assert RAM(16790) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16790))))  severity failure;
	assert RAM(16791) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(16791))))  severity failure;
	assert RAM(16792) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16792))))  severity failure;
	assert RAM(16793) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(16793))))  severity failure;
	assert RAM(16794) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16794))))  severity failure;
	assert RAM(16795) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16795))))  severity failure;
	assert RAM(16796) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16796))))  severity failure;
	assert RAM(16797) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16797))))  severity failure;
	assert RAM(16798) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16798))))  severity failure;
	assert RAM(16799) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16799))))  severity failure;
	assert RAM(16800) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16800))))  severity failure;
	assert RAM(16801) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16801))))  severity failure;
	assert RAM(16802) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16802))))  severity failure;
	assert RAM(16803) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(16803))))  severity failure;
	assert RAM(16804) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16804))))  severity failure;
	assert RAM(16805) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16805))))  severity failure;
	assert RAM(16806) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16806))))  severity failure;
	assert RAM(16807) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16807))))  severity failure;
	assert RAM(16808) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16808))))  severity failure;
	assert RAM(16809) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(16809))))  severity failure;
	assert RAM(16810) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(16810))))  severity failure;
	assert RAM(16811) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16811))))  severity failure;
	assert RAM(16812) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16812))))  severity failure;
	assert RAM(16813) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16813))))  severity failure;
	assert RAM(16814) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(16814))))  severity failure;
	assert RAM(16815) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16815))))  severity failure;
	assert RAM(16816) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16816))))  severity failure;
	assert RAM(16817) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16817))))  severity failure;
	assert RAM(16818) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(16818))))  severity failure;
	assert RAM(16819) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(16819))))  severity failure;
	assert RAM(16820) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16820))))  severity failure;
	assert RAM(16821) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16821))))  severity failure;
	assert RAM(16822) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(16822))))  severity failure;
	assert RAM(16823) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16823))))  severity failure;
	assert RAM(16824) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(16824))))  severity failure;
	assert RAM(16825) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(16825))))  severity failure;
	assert RAM(16826) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16826))))  severity failure;
	assert RAM(16827) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(16827))))  severity failure;
	assert RAM(16828) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16828))))  severity failure;
	assert RAM(16829) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16829))))  severity failure;
	assert RAM(16830) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16830))))  severity failure;
	assert RAM(16831) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16831))))  severity failure;
	assert RAM(16832) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16832))))  severity failure;
	assert RAM(16833) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16833))))  severity failure;
	assert RAM(16834) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16834))))  severity failure;
	assert RAM(16835) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16835))))  severity failure;
	assert RAM(16836) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16836))))  severity failure;
	assert RAM(16837) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16837))))  severity failure;
	assert RAM(16838) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16838))))  severity failure;
	assert RAM(16839) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16839))))  severity failure;
	assert RAM(16840) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(16840))))  severity failure;
	assert RAM(16841) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16841))))  severity failure;
	assert RAM(16842) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16842))))  severity failure;
	assert RAM(16843) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16843))))  severity failure;
	assert RAM(16844) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16844))))  severity failure;
	assert RAM(16845) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(16845))))  severity failure;
	assert RAM(16846) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(16846))))  severity failure;
	assert RAM(16847) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(16847))))  severity failure;
	assert RAM(16848) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16848))))  severity failure;
	assert RAM(16849) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16849))))  severity failure;
	assert RAM(16850) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16850))))  severity failure;
	assert RAM(16851) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16851))))  severity failure;
	assert RAM(16852) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16852))))  severity failure;
	assert RAM(16853) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16853))))  severity failure;
	assert RAM(16854) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16854))))  severity failure;
	assert RAM(16855) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16855))))  severity failure;
	assert RAM(16856) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(16856))))  severity failure;
	assert RAM(16857) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16857))))  severity failure;
	assert RAM(16858) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(16858))))  severity failure;
	assert RAM(16859) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16859))))  severity failure;
	assert RAM(16860) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16860))))  severity failure;
	assert RAM(16861) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(16861))))  severity failure;
	assert RAM(16862) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16862))))  severity failure;
	assert RAM(16863) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16863))))  severity failure;
	assert RAM(16864) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(16864))))  severity failure;
	assert RAM(16865) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16865))))  severity failure;
	assert RAM(16866) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16866))))  severity failure;
	assert RAM(16867) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16867))))  severity failure;
	assert RAM(16868) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16868))))  severity failure;
	assert RAM(16869) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16869))))  severity failure;
	assert RAM(16870) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(16870))))  severity failure;
	assert RAM(16871) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(16871))))  severity failure;
	assert RAM(16872) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16872))))  severity failure;
	assert RAM(16873) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16873))))  severity failure;
	assert RAM(16874) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16874))))  severity failure;
	assert RAM(16875) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16875))))  severity failure;
	assert RAM(16876) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16876))))  severity failure;
	assert RAM(16877) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(16877))))  severity failure;
	assert RAM(16878) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(16878))))  severity failure;
	assert RAM(16879) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(16879))))  severity failure;
	assert RAM(16880) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(16880))))  severity failure;
	assert RAM(16881) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16881))))  severity failure;
	assert RAM(16882) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16882))))  severity failure;
	assert RAM(16883) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(16883))))  severity failure;
	assert RAM(16884) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16884))))  severity failure;
	assert RAM(16885) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(16885))))  severity failure;
	assert RAM(16886) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(16886))))  severity failure;
	assert RAM(16887) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16887))))  severity failure;
	assert RAM(16888) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16888))))  severity failure;
	assert RAM(16889) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16889))))  severity failure;
	assert RAM(16890) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(16890))))  severity failure;
	assert RAM(16891) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(16891))))  severity failure;
	assert RAM(16892) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(16892))))  severity failure;
	assert RAM(16893) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16893))))  severity failure;
	assert RAM(16894) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16894))))  severity failure;
	assert RAM(16895) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16895))))  severity failure;
	assert RAM(16896) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16896))))  severity failure;
	assert RAM(16897) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16897))))  severity failure;
	assert RAM(16898) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16898))))  severity failure;
	assert RAM(16899) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16899))))  severity failure;
	assert RAM(16900) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16900))))  severity failure;
	assert RAM(16901) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(16901))))  severity failure;
	assert RAM(16902) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16902))))  severity failure;
	assert RAM(16903) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16903))))  severity failure;
	assert RAM(16904) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(16904))))  severity failure;
	assert RAM(16905) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(16905))))  severity failure;
	assert RAM(16906) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(16906))))  severity failure;
	assert RAM(16907) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(16907))))  severity failure;
	assert RAM(16908) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16908))))  severity failure;
	assert RAM(16909) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16909))))  severity failure;
	assert RAM(16910) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16910))))  severity failure;
	assert RAM(16911) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16911))))  severity failure;
	assert RAM(16912) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(16912))))  severity failure;
	assert RAM(16913) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16913))))  severity failure;
	assert RAM(16914) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16914))))  severity failure;
	assert RAM(16915) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(16915))))  severity failure;
	assert RAM(16916) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16916))))  severity failure;
	assert RAM(16917) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16917))))  severity failure;
	assert RAM(16918) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16918))))  severity failure;
	assert RAM(16919) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16919))))  severity failure;
	assert RAM(16920) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16920))))  severity failure;
	assert RAM(16921) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16921))))  severity failure;
	assert RAM(16922) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16922))))  severity failure;
	assert RAM(16923) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16923))))  severity failure;
	assert RAM(16924) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16924))))  severity failure;
	assert RAM(16925) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16925))))  severity failure;
	assert RAM(16926) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16926))))  severity failure;
	assert RAM(16927) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(16927))))  severity failure;
	assert RAM(16928) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16928))))  severity failure;
	assert RAM(16929) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(16929))))  severity failure;
	assert RAM(16930) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16930))))  severity failure;
	assert RAM(16931) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16931))))  severity failure;
	assert RAM(16932) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(16932))))  severity failure;
	assert RAM(16933) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16933))))  severity failure;
	assert RAM(16934) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(16934))))  severity failure;
	assert RAM(16935) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16935))))  severity failure;
	assert RAM(16936) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(16936))))  severity failure;
	assert RAM(16937) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16937))))  severity failure;
	assert RAM(16938) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(16938))))  severity failure;
	assert RAM(16939) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16939))))  severity failure;
	assert RAM(16940) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16940))))  severity failure;
	assert RAM(16941) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(16941))))  severity failure;
	assert RAM(16942) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16942))))  severity failure;
	assert RAM(16943) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16943))))  severity failure;
	assert RAM(16944) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16944))))  severity failure;
	assert RAM(16945) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16945))))  severity failure;
	assert RAM(16946) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16946))))  severity failure;
	assert RAM(16947) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(16947))))  severity failure;
	assert RAM(16948) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16948))))  severity failure;
	assert RAM(16949) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16949))))  severity failure;
	assert RAM(16950) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16950))))  severity failure;
	assert RAM(16951) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16951))))  severity failure;
	assert RAM(16952) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16952))))  severity failure;
	assert RAM(16953) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16953))))  severity failure;
	assert RAM(16954) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16954))))  severity failure;
	assert RAM(16955) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16955))))  severity failure;
	assert RAM(16956) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16956))))  severity failure;
	assert RAM(16957) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16957))))  severity failure;
	assert RAM(16958) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16958))))  severity failure;
	assert RAM(16959) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16959))))  severity failure;
	assert RAM(16960) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16960))))  severity failure;
	assert RAM(16961) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(16961))))  severity failure;
	assert RAM(16962) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16962))))  severity failure;
	assert RAM(16963) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16963))))  severity failure;
	assert RAM(16964) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16964))))  severity failure;
	assert RAM(16965) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(16965))))  severity failure;
	assert RAM(16966) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16966))))  severity failure;
	assert RAM(16967) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(16967))))  severity failure;
	assert RAM(16968) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16968))))  severity failure;
	assert RAM(16969) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(16969))))  severity failure;
	assert RAM(16970) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16970))))  severity failure;
	assert RAM(16971) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16971))))  severity failure;
	assert RAM(16972) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16972))))  severity failure;
	assert RAM(16973) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(16973))))  severity failure;
	assert RAM(16974) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(16974))))  severity failure;
	assert RAM(16975) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(16975))))  severity failure;
	assert RAM(16976) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16976))))  severity failure;
	assert RAM(16977) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16977))))  severity failure;
	assert RAM(16978) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16978))))  severity failure;
	assert RAM(16979) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16979))))  severity failure;
	assert RAM(16980) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(16980))))  severity failure;
	assert RAM(16981) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16981))))  severity failure;
	assert RAM(16982) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16982))))  severity failure;
	assert RAM(16983) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(16983))))  severity failure;
	assert RAM(16984) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16984))))  severity failure;
	assert RAM(16985) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16985))))  severity failure;
	assert RAM(16986) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16986))))  severity failure;
	assert RAM(16987) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16987))))  severity failure;
	assert RAM(16988) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16988))))  severity failure;
	assert RAM(16989) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16989))))  severity failure;
	assert RAM(16990) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16990))))  severity failure;
	assert RAM(16991) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16991))))  severity failure;
	assert RAM(16992) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(16992))))  severity failure;
	assert RAM(16993) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16993))))  severity failure;
	assert RAM(16994) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16994))))  severity failure;
	assert RAM(16995) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(16995))))  severity failure;
	assert RAM(16996) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16996))))  severity failure;
	assert RAM(16997) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16997))))  severity failure;
	assert RAM(16998) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16998))))  severity failure;
	assert RAM(16999) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16999))))  severity failure;
	assert RAM(17000) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17000))))  severity failure;
	assert RAM(17001) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17001))))  severity failure;
	assert RAM(17002) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17002))))  severity failure;
	assert RAM(17003) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17003))))  severity failure;
	assert RAM(17004) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17004))))  severity failure;
	assert RAM(17005) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17005))))  severity failure;
	assert RAM(17006) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17006))))  severity failure;
	assert RAM(17007) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(17007))))  severity failure;
	assert RAM(17008) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17008))))  severity failure;
	assert RAM(17009) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17009))))  severity failure;
	assert RAM(17010) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17010))))  severity failure;
	assert RAM(17011) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17011))))  severity failure;
	assert RAM(17012) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17012))))  severity failure;
	assert RAM(17013) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17013))))  severity failure;
	assert RAM(17014) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(17014))))  severity failure;
	assert RAM(17015) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(17015))))  severity failure;
	assert RAM(17016) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17016))))  severity failure;
	assert RAM(17017) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17017))))  severity failure;
	assert RAM(17018) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(17018))))  severity failure;
	assert RAM(17019) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17019))))  severity failure;
	assert RAM(17020) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17020))))  severity failure;
	assert RAM(17021) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(17021))))  severity failure;
	assert RAM(17022) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17022))))  severity failure;
	assert RAM(17023) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17023))))  severity failure;
	assert RAM(17024) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17024))))  severity failure;
	assert RAM(17025) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17025))))  severity failure;
	assert RAM(17026) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17026))))  severity failure;
	assert RAM(17027) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17027))))  severity failure;
	assert RAM(17028) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17028))))  severity failure;
	assert RAM(17029) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17029))))  severity failure;
	assert RAM(17030) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17030))))  severity failure;
	assert RAM(17031) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17031))))  severity failure;
	assert RAM(17032) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(17032))))  severity failure;
	assert RAM(17033) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17033))))  severity failure;
	assert RAM(17034) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17034))))  severity failure;
	assert RAM(17035) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17035))))  severity failure;
	assert RAM(17036) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17036))))  severity failure;
	assert RAM(17037) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17037))))  severity failure;
	assert RAM(17038) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17038))))  severity failure;
	assert RAM(17039) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17039))))  severity failure;
	assert RAM(17040) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17040))))  severity failure;
	assert RAM(17041) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17041))))  severity failure;
	assert RAM(17042) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(17042))))  severity failure;
	assert RAM(17043) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17043))))  severity failure;
	assert RAM(17044) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17044))))  severity failure;
	assert RAM(17045) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17045))))  severity failure;
	assert RAM(17046) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17046))))  severity failure;
	assert RAM(17047) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(17047))))  severity failure;
	assert RAM(17048) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(17048))))  severity failure;
	assert RAM(17049) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17049))))  severity failure;
	assert RAM(17050) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17050))))  severity failure;
	assert RAM(17051) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17051))))  severity failure;
	assert RAM(17052) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17052))))  severity failure;
	assert RAM(17053) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17053))))  severity failure;
	assert RAM(17054) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17054))))  severity failure;
	assert RAM(17055) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17055))))  severity failure;
	assert RAM(17056) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17056))))  severity failure;
	assert RAM(17057) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17057))))  severity failure;
	assert RAM(17058) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(17058))))  severity failure;
	assert RAM(17059) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17059))))  severity failure;
	assert RAM(17060) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17060))))  severity failure;
	assert RAM(17061) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17061))))  severity failure;
	assert RAM(17062) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17062))))  severity failure;
	assert RAM(17063) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(17063))))  severity failure;
	assert RAM(17064) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17064))))  severity failure;
	assert RAM(17065) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17065))))  severity failure;
	assert RAM(17066) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17066))))  severity failure;
	assert RAM(17067) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17067))))  severity failure;
	assert RAM(17068) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17068))))  severity failure;
	assert RAM(17069) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17069))))  severity failure;
	assert RAM(17070) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17070))))  severity failure;
	assert RAM(17071) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17071))))  severity failure;
	assert RAM(17072) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17072))))  severity failure;
	assert RAM(17073) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17073))))  severity failure;
	assert RAM(17074) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17074))))  severity failure;
	assert RAM(17075) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17075))))  severity failure;
	assert RAM(17076) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17076))))  severity failure;
	assert RAM(17077) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17077))))  severity failure;
	assert RAM(17078) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(17078))))  severity failure;
	assert RAM(17079) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17079))))  severity failure;
	assert RAM(17080) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17080))))  severity failure;
	assert RAM(17081) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(17081))))  severity failure;
	assert RAM(17082) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17082))))  severity failure;
	assert RAM(17083) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17083))))  severity failure;
	assert RAM(17084) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17084))))  severity failure;
	assert RAM(17085) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17085))))  severity failure;
	assert RAM(17086) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17086))))  severity failure;
	assert RAM(17087) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(17087))))  severity failure;
	assert RAM(17088) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17088))))  severity failure;
	assert RAM(17089) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17089))))  severity failure;
	assert RAM(17090) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17090))))  severity failure;
	assert RAM(17091) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17091))))  severity failure;
	assert RAM(17092) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17092))))  severity failure;
	assert RAM(17093) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17093))))  severity failure;
	assert RAM(17094) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17094))))  severity failure;
	assert RAM(17095) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17095))))  severity failure;
	assert RAM(17096) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17096))))  severity failure;
	assert RAM(17097) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17097))))  severity failure;
	assert RAM(17098) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17098))))  severity failure;
	assert RAM(17099) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17099))))  severity failure;
	assert RAM(17100) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17100))))  severity failure;
	assert RAM(17101) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17101))))  severity failure;
	assert RAM(17102) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17102))))  severity failure;
	assert RAM(17103) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17103))))  severity failure;
	assert RAM(17104) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17104))))  severity failure;
	assert RAM(17105) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17105))))  severity failure;
	assert RAM(17106) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17106))))  severity failure;
	assert RAM(17107) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17107))))  severity failure;
	assert RAM(17108) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17108))))  severity failure;
	assert RAM(17109) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17109))))  severity failure;
	assert RAM(17110) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(17110))))  severity failure;
	assert RAM(17111) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(17111))))  severity failure;
	assert RAM(17112) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17112))))  severity failure;
	assert RAM(17113) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17113))))  severity failure;
	assert RAM(17114) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17114))))  severity failure;
	assert RAM(17115) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17115))))  severity failure;
	assert RAM(17116) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17116))))  severity failure;
	assert RAM(17117) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17117))))  severity failure;
	assert RAM(17118) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17118))))  severity failure;
	assert RAM(17119) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17119))))  severity failure;
	assert RAM(17120) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17120))))  severity failure;
	assert RAM(17121) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17121))))  severity failure;
	assert RAM(17122) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17122))))  severity failure;
	assert RAM(17123) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17123))))  severity failure;
	assert RAM(17124) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17124))))  severity failure;
	assert RAM(17125) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(17125))))  severity failure;
	assert RAM(17126) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17126))))  severity failure;
	assert RAM(17127) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17127))))  severity failure;
	assert RAM(17128) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17128))))  severity failure;
	assert RAM(17129) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(17129))))  severity failure;
	assert RAM(17130) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17130))))  severity failure;
	assert RAM(17131) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(17131))))  severity failure;
	assert RAM(17132) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17132))))  severity failure;
	assert RAM(17133) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17133))))  severity failure;
	assert RAM(17134) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17134))))  severity failure;
	assert RAM(17135) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17135))))  severity failure;
	assert RAM(17136) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17136))))  severity failure;
	assert RAM(17137) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17137))))  severity failure;
	assert RAM(17138) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(17138))))  severity failure;
	assert RAM(17139) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17139))))  severity failure;
	assert RAM(17140) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17140))))  severity failure;
	assert RAM(17141) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17141))))  severity failure;
	assert RAM(17142) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17142))))  severity failure;
	assert RAM(17143) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17143))))  severity failure;
	assert RAM(17144) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17144))))  severity failure;
	assert RAM(17145) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17145))))  severity failure;
	assert RAM(17146) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17146))))  severity failure;
	assert RAM(17147) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17147))))  severity failure;
	assert RAM(17148) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17148))))  severity failure;
	assert RAM(17149) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17149))))  severity failure;
	assert RAM(17150) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17150))))  severity failure;
	assert RAM(17151) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17151))))  severity failure;
	assert RAM(17152) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17152))))  severity failure;
	assert RAM(17153) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17153))))  severity failure;
	assert RAM(17154) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17154))))  severity failure;
	assert RAM(17155) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17155))))  severity failure;
	assert RAM(17156) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17156))))  severity failure;
	assert RAM(17157) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17157))))  severity failure;
	assert RAM(17158) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17158))))  severity failure;
	assert RAM(17159) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17159))))  severity failure;
	assert RAM(17160) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17160))))  severity failure;
	assert RAM(17161) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17161))))  severity failure;
	assert RAM(17162) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17162))))  severity failure;
	assert RAM(17163) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17163))))  severity failure;
	assert RAM(17164) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17164))))  severity failure;
	assert RAM(17165) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17165))))  severity failure;
	assert RAM(17166) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17166))))  severity failure;
	assert RAM(17167) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17167))))  severity failure;
	assert RAM(17168) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(17168))))  severity failure;
	assert RAM(17169) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17169))))  severity failure;
	assert RAM(17170) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(17170))))  severity failure;
	assert RAM(17171) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17171))))  severity failure;
	assert RAM(17172) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17172))))  severity failure;
	assert RAM(17173) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17173))))  severity failure;
	assert RAM(17174) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17174))))  severity failure;
	assert RAM(17175) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17175))))  severity failure;
	assert RAM(17176) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17176))))  severity failure;
	assert RAM(17177) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17177))))  severity failure;
	assert RAM(17178) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17178))))  severity failure;
	assert RAM(17179) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17179))))  severity failure;
	assert RAM(17180) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17180))))  severity failure;
	assert RAM(17181) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17181))))  severity failure;
	assert RAM(17182) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17182))))  severity failure;
	assert RAM(17183) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17183))))  severity failure;
	assert RAM(17184) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17184))))  severity failure;
	assert RAM(17185) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17185))))  severity failure;
	assert RAM(17186) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17186))))  severity failure;
	assert RAM(17187) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17187))))  severity failure;
	assert RAM(17188) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17188))))  severity failure;
	assert RAM(17189) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(17189))))  severity failure;
	assert RAM(17190) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(17190))))  severity failure;
	assert RAM(17191) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17191))))  severity failure;
	assert RAM(17192) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17192))))  severity failure;
	assert RAM(17193) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17193))))  severity failure;
	assert RAM(17194) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17194))))  severity failure;
	assert RAM(17195) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17195))))  severity failure;
	assert RAM(17196) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17196))))  severity failure;
	assert RAM(17197) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17197))))  severity failure;
	assert RAM(17198) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17198))))  severity failure;
	assert RAM(17199) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17199))))  severity failure;
	assert RAM(17200) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17200))))  severity failure;
	assert RAM(17201) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(17201))))  severity failure;
	assert RAM(17202) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17202))))  severity failure;
	assert RAM(17203) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17203))))  severity failure;
	assert RAM(17204) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17204))))  severity failure;
	assert RAM(17205) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(17205))))  severity failure;
	assert RAM(17206) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17206))))  severity failure;
	assert RAM(17207) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17207))))  severity failure;
	assert RAM(17208) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17208))))  severity failure;
	assert RAM(17209) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(17209))))  severity failure;
	assert RAM(17210) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17210))))  severity failure;
	assert RAM(17211) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17211))))  severity failure;
	assert RAM(17212) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(17212))))  severity failure;
	assert RAM(17213) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17213))))  severity failure;
	assert RAM(17214) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17214))))  severity failure;
	assert RAM(17215) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17215))))  severity failure;
	assert RAM(17216) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17216))))  severity failure;
	assert RAM(17217) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17217))))  severity failure;
	assert RAM(17218) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17218))))  severity failure;
	assert RAM(17219) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17219))))  severity failure;
	assert RAM(17220) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17220))))  severity failure;
	assert RAM(17221) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17221))))  severity failure;
	assert RAM(17222) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(17222))))  severity failure;
	assert RAM(17223) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17223))))  severity failure;
	assert RAM(17224) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(17224))))  severity failure;
	assert RAM(17225) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17225))))  severity failure;
	assert RAM(17226) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17226))))  severity failure;
	assert RAM(17227) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17227))))  severity failure;
	assert RAM(17228) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17228))))  severity failure;
	assert RAM(17229) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17229))))  severity failure;
	assert RAM(17230) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17230))))  severity failure;
	assert RAM(17231) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17231))))  severity failure;
	assert RAM(17232) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17232))))  severity failure;
	assert RAM(17233) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17233))))  severity failure;
	assert RAM(17234) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17234))))  severity failure;
	assert RAM(17235) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17235))))  severity failure;
	assert RAM(17236) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17236))))  severity failure;
	assert RAM(17237) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17237))))  severity failure;
	assert RAM(17238) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17238))))  severity failure;
	assert RAM(17239) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17239))))  severity failure;
	assert RAM(17240) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17240))))  severity failure;
	assert RAM(17241) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17241))))  severity failure;
	assert RAM(17242) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17242))))  severity failure;
	assert RAM(17243) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17243))))  severity failure;
	assert RAM(17244) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(17244))))  severity failure;
	assert RAM(17245) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17245))))  severity failure;
	assert RAM(17246) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17246))))  severity failure;
	assert RAM(17247) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17247))))  severity failure;
	assert RAM(17248) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17248))))  severity failure;
	assert RAM(17249) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(17249))))  severity failure;
	assert RAM(17250) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17250))))  severity failure;
	assert RAM(17251) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17251))))  severity failure;
	assert RAM(17252) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17252))))  severity failure;
	assert RAM(17253) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(17253))))  severity failure;
	assert RAM(17254) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17254))))  severity failure;
	assert RAM(17255) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17255))))  severity failure;
	assert RAM(17256) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17256))))  severity failure;
	assert RAM(17257) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17257))))  severity failure;
	assert RAM(17258) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17258))))  severity failure;
	assert RAM(17259) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17259))))  severity failure;
	assert RAM(17260) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17260))))  severity failure;
	assert RAM(17261) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17261))))  severity failure;
	assert RAM(17262) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(17262))))  severity failure;
	assert RAM(17263) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17263))))  severity failure;
	assert RAM(17264) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17264))))  severity failure;
	assert RAM(17265) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17265))))  severity failure;
	assert RAM(17266) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17266))))  severity failure;
	assert RAM(17267) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17267))))  severity failure;
	assert RAM(17268) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17268))))  severity failure;
	assert RAM(17269) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17269))))  severity failure;
	assert RAM(17270) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17270))))  severity failure;
	assert RAM(17271) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(17271))))  severity failure;
	assert RAM(17272) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(17272))))  severity failure;
	assert RAM(17273) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17273))))  severity failure;
	assert RAM(17274) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17274))))  severity failure;
	assert RAM(17275) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17275))))  severity failure;
	assert RAM(17276) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17276))))  severity failure;
	assert RAM(17277) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17277))))  severity failure;
	assert RAM(17278) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17278))))  severity failure;
	assert RAM(17279) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17279))))  severity failure;
	assert RAM(17280) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17280))))  severity failure;
	assert RAM(17281) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17281))))  severity failure;
	assert RAM(17282) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17282))))  severity failure;
	assert RAM(17283) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17283))))  severity failure;
	assert RAM(17284) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17284))))  severity failure;
	assert RAM(17285) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17285))))  severity failure;
	assert RAM(17286) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17286))))  severity failure;
	assert RAM(17287) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17287))))  severity failure;
	assert RAM(17288) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17288))))  severity failure;
	assert RAM(17289) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17289))))  severity failure;
	assert RAM(17290) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17290))))  severity failure;
	assert RAM(17291) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17291))))  severity failure;
	assert RAM(17292) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17292))))  severity failure;
	assert RAM(17293) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17293))))  severity failure;
	assert RAM(17294) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17294))))  severity failure;
	assert RAM(17295) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17295))))  severity failure;
	assert RAM(17296) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17296))))  severity failure;
	assert RAM(17297) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17297))))  severity failure;
	assert RAM(17298) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17298))))  severity failure;
	assert RAM(17299) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17299))))  severity failure;
	assert RAM(17300) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17300))))  severity failure;
	assert RAM(17301) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17301))))  severity failure;
	assert RAM(17302) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17302))))  severity failure;
	assert RAM(17303) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17303))))  severity failure;
	assert RAM(17304) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17304))))  severity failure;
	assert RAM(17305) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17305))))  severity failure;
	assert RAM(17306) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17306))))  severity failure;
	assert RAM(17307) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17307))))  severity failure;
	assert RAM(17308) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17308))))  severity failure;
	assert RAM(17309) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(17309))))  severity failure;
	assert RAM(17310) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17310))))  severity failure;
	assert RAM(17311) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17311))))  severity failure;
	assert RAM(17312) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17312))))  severity failure;
	assert RAM(17313) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17313))))  severity failure;
	assert RAM(17314) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17314))))  severity failure;
	assert RAM(17315) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17315))))  severity failure;
	assert RAM(17316) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17316))))  severity failure;
	assert RAM(17317) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(17317))))  severity failure;
	assert RAM(17318) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17318))))  severity failure;
	assert RAM(17319) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17319))))  severity failure;
	assert RAM(17320) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(17320))))  severity failure;
	assert RAM(17321) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17321))))  severity failure;
	assert RAM(17322) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(17322))))  severity failure;
	assert RAM(17323) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17323))))  severity failure;
	assert RAM(17324) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17324))))  severity failure;
	assert RAM(17325) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17325))))  severity failure;
	assert RAM(17326) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17326))))  severity failure;
	assert RAM(17327) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17327))))  severity failure;
	assert RAM(17328) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17328))))  severity failure;
	assert RAM(17329) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17329))))  severity failure;
	assert RAM(17330) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17330))))  severity failure;
	assert RAM(17331) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17331))))  severity failure;
	assert RAM(17332) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17332))))  severity failure;
	assert RAM(17333) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17333))))  severity failure;
	assert RAM(17334) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17334))))  severity failure;
	assert RAM(17335) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17335))))  severity failure;
	assert RAM(17336) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17336))))  severity failure;
	assert RAM(17337) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17337))))  severity failure;
	assert RAM(17338) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17338))))  severity failure;
	assert RAM(17339) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17339))))  severity failure;
	assert RAM(17340) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17340))))  severity failure;
	assert RAM(17341) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17341))))  severity failure;
	assert RAM(17342) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(17342))))  severity failure;
	assert RAM(17343) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17343))))  severity failure;
	assert RAM(17344) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17344))))  severity failure;
	assert RAM(17345) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17345))))  severity failure;
	assert RAM(17346) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17346))))  severity failure;
	assert RAM(17347) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17347))))  severity failure;
	assert RAM(17348) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17348))))  severity failure;
	assert RAM(17349) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17349))))  severity failure;
	assert RAM(17350) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17350))))  severity failure;
	assert RAM(17351) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17351))))  severity failure;
	assert RAM(17352) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17352))))  severity failure;
	assert RAM(17353) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17353))))  severity failure;
	assert RAM(17354) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17354))))  severity failure;
	assert RAM(17355) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(17355))))  severity failure;
	assert RAM(17356) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17356))))  severity failure;
	assert RAM(17357) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17357))))  severity failure;
	assert RAM(17358) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17358))))  severity failure;
	assert RAM(17359) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17359))))  severity failure;
	assert RAM(17360) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17360))))  severity failure;
	assert RAM(17361) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17361))))  severity failure;
	assert RAM(17362) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17362))))  severity failure;
	assert RAM(17363) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17363))))  severity failure;
	assert RAM(17364) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17364))))  severity failure;
	assert RAM(17365) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17365))))  severity failure;
	assert RAM(17366) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17366))))  severity failure;
	assert RAM(17367) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17367))))  severity failure;
	assert RAM(17368) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17368))))  severity failure;
	assert RAM(17369) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17369))))  severity failure;
	assert RAM(17370) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17370))))  severity failure;
	assert RAM(17371) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17371))))  severity failure;
	assert RAM(17372) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17372))))  severity failure;
	assert RAM(17373) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17373))))  severity failure;
	assert RAM(17374) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(17374))))  severity failure;
	assert RAM(17375) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17375))))  severity failure;
	assert RAM(17376) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17376))))  severity failure;
	assert RAM(17377) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(17377))))  severity failure;
	assert RAM(17378) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(17378))))  severity failure;
	assert RAM(17379) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17379))))  severity failure;
	assert RAM(17380) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17380))))  severity failure;
	assert RAM(17381) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17381))))  severity failure;
	assert RAM(17382) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17382))))  severity failure;
	assert RAM(17383) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17383))))  severity failure;
	assert RAM(17384) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17384))))  severity failure;
	assert RAM(17385) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17385))))  severity failure;
	assert RAM(17386) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17386))))  severity failure;
	assert RAM(17387) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17387))))  severity failure;
	assert RAM(17388) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17388))))  severity failure;
	assert RAM(17389) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17389))))  severity failure;
	assert RAM(17390) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17390))))  severity failure;
	assert RAM(17391) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17391))))  severity failure;
	assert RAM(17392) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17392))))  severity failure;
	assert RAM(17393) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17393))))  severity failure;
	assert RAM(17394) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17394))))  severity failure;
	assert RAM(17395) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17395))))  severity failure;
	assert RAM(17396) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17396))))  severity failure;
	assert RAM(17397) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17397))))  severity failure;
	assert RAM(17398) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17398))))  severity failure;
	assert RAM(17399) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17399))))  severity failure;
	assert RAM(17400) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17400))))  severity failure;
	assert RAM(17401) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17401))))  severity failure;
	assert RAM(17402) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17402))))  severity failure;
	assert RAM(17403) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17403))))  severity failure;
	assert RAM(17404) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17404))))  severity failure;
	assert RAM(17405) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17405))))  severity failure;
	assert RAM(17406) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17406))))  severity failure;
	assert RAM(17407) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17407))))  severity failure;
	assert RAM(17408) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17408))))  severity failure;
	assert RAM(17409) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17409))))  severity failure;
	assert RAM(17410) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(17410))))  severity failure;
	assert RAM(17411) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17411))))  severity failure;
	assert RAM(17412) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(17412))))  severity failure;
	assert RAM(17413) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17413))))  severity failure;
	assert RAM(17414) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17414))))  severity failure;
	assert RAM(17415) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17415))))  severity failure;
	assert RAM(17416) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17416))))  severity failure;
	assert RAM(17417) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17417))))  severity failure;
	assert RAM(17418) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17418))))  severity failure;
	assert RAM(17419) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(17419))))  severity failure;
	assert RAM(17420) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17420))))  severity failure;
	assert RAM(17421) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17421))))  severity failure;
	assert RAM(17422) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17422))))  severity failure;
	assert RAM(17423) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17423))))  severity failure;
	assert RAM(17424) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(17424))))  severity failure;
	assert RAM(17425) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17425))))  severity failure;
	assert RAM(17426) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17426))))  severity failure;
	assert RAM(17427) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17427))))  severity failure;
	assert RAM(17428) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17428))))  severity failure;
	assert RAM(17429) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17429))))  severity failure;
	assert RAM(17430) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17430))))  severity failure;
	assert RAM(17431) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17431))))  severity failure;
	assert RAM(17432) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(17432))))  severity failure;
	assert RAM(17433) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17433))))  severity failure;
	assert RAM(17434) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17434))))  severity failure;
	assert RAM(17435) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17435))))  severity failure;
	assert RAM(17436) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17436))))  severity failure;
	assert RAM(17437) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17437))))  severity failure;
	assert RAM(17438) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17438))))  severity failure;
	assert RAM(17439) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(17439))))  severity failure;
	assert RAM(17440) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17440))))  severity failure;
	assert RAM(17441) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17441))))  severity failure;
	assert RAM(17442) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17442))))  severity failure;
	assert RAM(17443) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(17443))))  severity failure;
	assert RAM(17444) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17444))))  severity failure;
	assert RAM(17445) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17445))))  severity failure;
	assert RAM(17446) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17446))))  severity failure;
	assert RAM(17447) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17447))))  severity failure;
	assert RAM(17448) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17448))))  severity failure;
	assert RAM(17449) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17449))))  severity failure;
	assert RAM(17450) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(17450))))  severity failure;
	assert RAM(17451) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17451))))  severity failure;
	assert RAM(17452) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17452))))  severity failure;
	assert RAM(17453) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(17453))))  severity failure;
	assert RAM(17454) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17454))))  severity failure;
	assert RAM(17455) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17455))))  severity failure;
	assert RAM(17456) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17456))))  severity failure;
	assert RAM(17457) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17457))))  severity failure;
	assert RAM(17458) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17458))))  severity failure;
	assert RAM(17459) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17459))))  severity failure;
	assert RAM(17460) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(17460))))  severity failure;
	assert RAM(17461) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17461))))  severity failure;
	assert RAM(17462) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17462))))  severity failure;
	assert RAM(17463) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17463))))  severity failure;
	assert RAM(17464) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17464))))  severity failure;
	assert RAM(17465) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17465))))  severity failure;
	assert RAM(17466) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(17466))))  severity failure;
	assert RAM(17467) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17467))))  severity failure;
	assert RAM(17468) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17468))))  severity failure;
	assert RAM(17469) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17469))))  severity failure;
	assert RAM(17470) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17470))))  severity failure;
	assert RAM(17471) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17471))))  severity failure;
	assert RAM(17472) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17472))))  severity failure;
	assert RAM(17473) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17473))))  severity failure;
	assert RAM(17474) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17474))))  severity failure;
	assert RAM(17475) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17475))))  severity failure;
	assert RAM(17476) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17476))))  severity failure;
	assert RAM(17477) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17477))))  severity failure;
	assert RAM(17478) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17478))))  severity failure;
	assert RAM(17479) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17479))))  severity failure;
	assert RAM(17480) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17480))))  severity failure;
	assert RAM(17481) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17481))))  severity failure;
	assert RAM(17482) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17482))))  severity failure;
	assert RAM(17483) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17483))))  severity failure;
	assert RAM(17484) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(17484))))  severity failure;
	assert RAM(17485) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(17485))))  severity failure;
	assert RAM(17486) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17486))))  severity failure;
	assert RAM(17487) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(17487))))  severity failure;
	assert RAM(17488) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17488))))  severity failure;
	assert RAM(17489) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17489))))  severity failure;
	assert RAM(17490) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17490))))  severity failure;
	assert RAM(17491) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17491))))  severity failure;
	assert RAM(17492) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(17492))))  severity failure;
	assert RAM(17493) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17493))))  severity failure;
	assert RAM(17494) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17494))))  severity failure;
	assert RAM(17495) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17495))))  severity failure;
	assert RAM(17496) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17496))))  severity failure;
	assert RAM(17497) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17497))))  severity failure;
	assert RAM(17498) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17498))))  severity failure;
	assert RAM(17499) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17499))))  severity failure;
	assert RAM(17500) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17500))))  severity failure;
	assert RAM(17501) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17501))))  severity failure;
	assert RAM(17502) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(17502))))  severity failure;
	assert RAM(17503) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17503))))  severity failure;
	assert RAM(17504) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17504))))  severity failure;
	assert RAM(17505) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17505))))  severity failure;
	assert RAM(17506) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17506))))  severity failure;
	assert RAM(17507) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17507))))  severity failure;
	assert RAM(17508) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17508))))  severity failure;
	assert RAM(17509) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17509))))  severity failure;
	assert RAM(17510) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17510))))  severity failure;
	assert RAM(17511) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17511))))  severity failure;
	assert RAM(17512) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17512))))  severity failure;
	assert RAM(17513) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17513))))  severity failure;
	assert RAM(17514) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17514))))  severity failure;
	assert RAM(17515) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17515))))  severity failure;
	assert RAM(17516) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17516))))  severity failure;
	assert RAM(17517) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17517))))  severity failure;
	assert RAM(17518) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17518))))  severity failure;
	assert RAM(17519) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17519))))  severity failure;
	assert RAM(17520) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17520))))  severity failure;
	assert RAM(17521) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17521))))  severity failure;
	assert RAM(17522) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(17522))))  severity failure;
	assert RAM(17523) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17523))))  severity failure;
	assert RAM(17524) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17524))))  severity failure;
	assert RAM(17525) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17525))))  severity failure;
	assert RAM(17526) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17526))))  severity failure;
	assert RAM(17527) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17527))))  severity failure;
	assert RAM(17528) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17528))))  severity failure;
	assert RAM(17529) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17529))))  severity failure;
	assert RAM(17530) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17530))))  severity failure;
	assert RAM(17531) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17531))))  severity failure;
	assert RAM(17532) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17532))))  severity failure;
	assert RAM(17533) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17533))))  severity failure;
	assert RAM(17534) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17534))))  severity failure;
	assert RAM(17535) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17535))))  severity failure;
	assert RAM(17536) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17536))))  severity failure;
	assert RAM(17537) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17537))))  severity failure;
	assert RAM(17538) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(17538))))  severity failure;
	assert RAM(17539) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17539))))  severity failure;
	assert RAM(17540) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17540))))  severity failure;
	assert RAM(17541) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17541))))  severity failure;
	assert RAM(17542) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17542))))  severity failure;
	assert RAM(17543) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17543))))  severity failure;
	assert RAM(17544) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17544))))  severity failure;
	assert RAM(17545) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17545))))  severity failure;
	assert RAM(17546) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17546))))  severity failure;
	assert RAM(17547) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17547))))  severity failure;
	assert RAM(17548) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17548))))  severity failure;
	assert RAM(17549) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17549))))  severity failure;
	assert RAM(17550) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17550))))  severity failure;
	assert RAM(17551) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(17551))))  severity failure;
	assert RAM(17552) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(17552))))  severity failure;
	assert RAM(17553) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17553))))  severity failure;
	assert RAM(17554) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(17554))))  severity failure;
	assert RAM(17555) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17555))))  severity failure;
	assert RAM(17556) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17556))))  severity failure;
	assert RAM(17557) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17557))))  severity failure;
	assert RAM(17558) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17558))))  severity failure;
	assert RAM(17559) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17559))))  severity failure;
	assert RAM(17560) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17560))))  severity failure;
	assert RAM(17561) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17561))))  severity failure;
	assert RAM(17562) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(17562))))  severity failure;
	assert RAM(17563) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(17563))))  severity failure;
	assert RAM(17564) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17564))))  severity failure;
	assert RAM(17565) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17565))))  severity failure;
	assert RAM(17566) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17566))))  severity failure;
	assert RAM(17567) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17567))))  severity failure;
	assert RAM(17568) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(17568))))  severity failure;
	assert RAM(17569) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17569))))  severity failure;
	assert RAM(17570) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17570))))  severity failure;
	assert RAM(17571) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17571))))  severity failure;
	assert RAM(17572) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(17572))))  severity failure;
	assert RAM(17573) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17573))))  severity failure;
	assert RAM(17574) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17574))))  severity failure;
	assert RAM(17575) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17575))))  severity failure;
	assert RAM(17576) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17576))))  severity failure;
	assert RAM(17577) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17577))))  severity failure;
	assert RAM(17578) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17578))))  severity failure;
	assert RAM(17579) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(17579))))  severity failure;
	assert RAM(17580) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17580))))  severity failure;
	assert RAM(17581) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17581))))  severity failure;
	assert RAM(17582) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(17582))))  severity failure;
	assert RAM(17583) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17583))))  severity failure;
	assert RAM(17584) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17584))))  severity failure;
	assert RAM(17585) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17585))))  severity failure;
	assert RAM(17586) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17586))))  severity failure;
	assert RAM(17587) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17587))))  severity failure;
	assert RAM(17588) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17588))))  severity failure;
	assert RAM(17589) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17589))))  severity failure;
	assert RAM(17590) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17590))))  severity failure;
	assert RAM(17591) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17591))))  severity failure;
	assert RAM(17592) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17592))))  severity failure;
	assert RAM(17593) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17593))))  severity failure;
	assert RAM(17594) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17594))))  severity failure;
	assert RAM(17595) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17595))))  severity failure;
	assert RAM(17596) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17596))))  severity failure;
	assert RAM(17597) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17597))))  severity failure;
	assert RAM(17598) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17598))))  severity failure;
	assert RAM(17599) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17599))))  severity failure;
	assert RAM(17600) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17600))))  severity failure;
	assert RAM(17601) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17601))))  severity failure;
	assert RAM(17602) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17602))))  severity failure;
	assert RAM(17603) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17603))))  severity failure;
	assert RAM(17604) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(17604))))  severity failure;
	assert RAM(17605) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17605))))  severity failure;
	assert RAM(17606) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17606))))  severity failure;
	assert RAM(17607) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17607))))  severity failure;
	assert RAM(17608) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17608))))  severity failure;
	assert RAM(17609) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17609))))  severity failure;
	assert RAM(17610) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17610))))  severity failure;
	assert RAM(17611) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17611))))  severity failure;
	assert RAM(17612) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17612))))  severity failure;
	assert RAM(17613) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(17613))))  severity failure;
	assert RAM(17614) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17614))))  severity failure;
	assert RAM(17615) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17615))))  severity failure;
	assert RAM(17616) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17616))))  severity failure;
	assert RAM(17617) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17617))))  severity failure;
	assert RAM(17618) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17618))))  severity failure;
	assert RAM(17619) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17619))))  severity failure;
	assert RAM(17620) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17620))))  severity failure;
	assert RAM(17621) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17621))))  severity failure;
	assert RAM(17622) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(17622))))  severity failure;
	assert RAM(17623) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17623))))  severity failure;
	assert RAM(17624) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17624))))  severity failure;
	assert RAM(17625) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17625))))  severity failure;
	assert RAM(17626) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17626))))  severity failure;
	assert RAM(17627) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17627))))  severity failure;
	assert RAM(17628) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(17628))))  severity failure;
	assert RAM(17629) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17629))))  severity failure;
	assert RAM(17630) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17630))))  severity failure;
	assert RAM(17631) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17631))))  severity failure;
	assert RAM(17632) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17632))))  severity failure;
	assert RAM(17633) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17633))))  severity failure;
	assert RAM(17634) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(17634))))  severity failure;
	assert RAM(17635) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(17635))))  severity failure;
	assert RAM(17636) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17636))))  severity failure;
	assert RAM(17637) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17637))))  severity failure;
	assert RAM(17638) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17638))))  severity failure;
	assert RAM(17639) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17639))))  severity failure;
	assert RAM(17640) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17640))))  severity failure;
	assert RAM(17641) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17641))))  severity failure;
	assert RAM(17642) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17642))))  severity failure;
	assert RAM(17643) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17643))))  severity failure;
	assert RAM(17644) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17644))))  severity failure;
	assert RAM(17645) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17645))))  severity failure;
	assert RAM(17646) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17646))))  severity failure;
	assert RAM(17647) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17647))))  severity failure;
	assert RAM(17648) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(17648))))  severity failure;
	assert RAM(17649) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17649))))  severity failure;
	assert RAM(17650) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17650))))  severity failure;
	assert RAM(17651) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17651))))  severity failure;
	assert RAM(17652) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(17652))))  severity failure;
	assert RAM(17653) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17653))))  severity failure;
	assert RAM(17654) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17654))))  severity failure;
	assert RAM(17655) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17655))))  severity failure;
	assert RAM(17656) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17656))))  severity failure;
	assert RAM(17657) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17657))))  severity failure;
	assert RAM(17658) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17658))))  severity failure;
	assert RAM(17659) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17659))))  severity failure;
	assert RAM(17660) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17660))))  severity failure;
	assert RAM(17661) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17661))))  severity failure;
	assert RAM(17662) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17662))))  severity failure;
	assert RAM(17663) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17663))))  severity failure;
	assert RAM(17664) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17664))))  severity failure;
	assert RAM(17665) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17665))))  severity failure;
	assert RAM(17666) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17666))))  severity failure;
	assert RAM(17667) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17667))))  severity failure;
	assert RAM(17668) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17668))))  severity failure;
	assert RAM(17669) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17669))))  severity failure;
	assert RAM(17670) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17670))))  severity failure;
	assert RAM(17671) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17671))))  severity failure;
	assert RAM(17672) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(17672))))  severity failure;
	assert RAM(17673) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17673))))  severity failure;
	assert RAM(17674) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17674))))  severity failure;
	assert RAM(17675) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(17675))))  severity failure;
	assert RAM(17676) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(17676))))  severity failure;
	assert RAM(17677) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17677))))  severity failure;
	assert RAM(17678) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17678))))  severity failure;
	assert RAM(17679) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17679))))  severity failure;
	assert RAM(17680) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17680))))  severity failure;
	assert RAM(17681) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17681))))  severity failure;
	assert RAM(17682) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17682))))  severity failure;
	assert RAM(17683) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17683))))  severity failure;
	assert RAM(17684) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(17684))))  severity failure;
	assert RAM(17685) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17685))))  severity failure;
	assert RAM(17686) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(17686))))  severity failure;
	assert RAM(17687) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17687))))  severity failure;
	assert RAM(17688) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17688))))  severity failure;
	assert RAM(17689) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17689))))  severity failure;
	assert RAM(17690) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17690))))  severity failure;
	assert RAM(17691) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17691))))  severity failure;
	assert RAM(17692) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17692))))  severity failure;
	assert RAM(17693) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17693))))  severity failure;
	assert RAM(17694) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17694))))  severity failure;
	assert RAM(17695) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17695))))  severity failure;
	assert RAM(17696) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(17696))))  severity failure;
	assert RAM(17697) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17697))))  severity failure;
	assert RAM(17698) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17698))))  severity failure;
	assert RAM(17699) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17699))))  severity failure;
	assert RAM(17700) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17700))))  severity failure;
	assert RAM(17701) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17701))))  severity failure;
	assert RAM(17702) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(17702))))  severity failure;
	assert RAM(17703) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17703))))  severity failure;
	assert RAM(17704) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17704))))  severity failure;
	assert RAM(17705) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17705))))  severity failure;
	assert RAM(17706) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17706))))  severity failure;
	assert RAM(17707) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17707))))  severity failure;
	assert RAM(17708) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(17708))))  severity failure;
	assert RAM(17709) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(17709))))  severity failure;
	assert RAM(17710) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17710))))  severity failure;
	assert RAM(17711) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17711))))  severity failure;
	assert RAM(17712) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17712))))  severity failure;
	assert RAM(17713) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17713))))  severity failure;
	assert RAM(17714) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17714))))  severity failure;
	assert RAM(17715) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17715))))  severity failure;
	assert RAM(17716) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17716))))  severity failure;
	assert RAM(17717) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17717))))  severity failure;
	assert RAM(17718) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17718))))  severity failure;
	assert RAM(17719) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17719))))  severity failure;
	assert RAM(17720) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17720))))  severity failure;
	assert RAM(17721) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17721))))  severity failure;
	assert RAM(17722) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17722))))  severity failure;
	assert RAM(17723) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17723))))  severity failure;
	assert RAM(17724) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17724))))  severity failure;
	assert RAM(17725) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17725))))  severity failure;
	assert RAM(17726) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17726))))  severity failure;
	assert RAM(17727) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17727))))  severity failure;
	assert RAM(17728) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17728))))  severity failure;
	assert RAM(17729) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17729))))  severity failure;
	assert RAM(17730) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17730))))  severity failure;
	assert RAM(17731) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17731))))  severity failure;
	assert RAM(17732) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17732))))  severity failure;
	assert RAM(17733) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17733))))  severity failure;
	assert RAM(17734) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17734))))  severity failure;
	assert RAM(17735) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17735))))  severity failure;
	assert RAM(17736) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17736))))  severity failure;
	assert RAM(17737) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17737))))  severity failure;
	assert RAM(17738) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17738))))  severity failure;
	assert RAM(17739) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17739))))  severity failure;
	assert RAM(17740) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17740))))  severity failure;
	assert RAM(17741) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17741))))  severity failure;
	assert RAM(17742) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17742))))  severity failure;
	assert RAM(17743) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17743))))  severity failure;
	assert RAM(17744) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(17744))))  severity failure;
	assert RAM(17745) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17745))))  severity failure;
	assert RAM(17746) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17746))))  severity failure;
	assert RAM(17747) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17747))))  severity failure;
	assert RAM(17748) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17748))))  severity failure;
	assert RAM(17749) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17749))))  severity failure;
	assert RAM(17750) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17750))))  severity failure;
	assert RAM(17751) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17751))))  severity failure;
	assert RAM(17752) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17752))))  severity failure;
	assert RAM(17753) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17753))))  severity failure;
	assert RAM(17754) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17754))))  severity failure;
	assert RAM(17755) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17755))))  severity failure;
	assert RAM(17756) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17756))))  severity failure;
	assert RAM(17757) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17757))))  severity failure;
	assert RAM(17758) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17758))))  severity failure;
	assert RAM(17759) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17759))))  severity failure;
	assert RAM(17760) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17760))))  severity failure;
	assert RAM(17761) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17761))))  severity failure;
	assert RAM(17762) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(17762))))  severity failure;
	assert RAM(17763) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17763))))  severity failure;
	assert RAM(17764) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17764))))  severity failure;
	assert RAM(17765) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17765))))  severity failure;
	assert RAM(17766) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17766))))  severity failure;
	assert RAM(17767) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17767))))  severity failure;
	assert RAM(17768) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(17768))))  severity failure;
	assert RAM(17769) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17769))))  severity failure;
	assert RAM(17770) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17770))))  severity failure;
	assert RAM(17771) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17771))))  severity failure;
	assert RAM(17772) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17772))))  severity failure;
	assert RAM(17773) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17773))))  severity failure;
	assert RAM(17774) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17774))))  severity failure;
	assert RAM(17775) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17775))))  severity failure;
	assert RAM(17776) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(17776))))  severity failure;
	assert RAM(17777) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(17777))))  severity failure;
	assert RAM(17778) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17778))))  severity failure;
	assert RAM(17779) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17779))))  severity failure;
	assert RAM(17780) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17780))))  severity failure;
	assert RAM(17781) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17781))))  severity failure;
	assert RAM(17782) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17782))))  severity failure;
	assert RAM(17783) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17783))))  severity failure;
	assert RAM(17784) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17784))))  severity failure;
	assert RAM(17785) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17785))))  severity failure;
	assert RAM(17786) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17786))))  severity failure;
	assert RAM(17787) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17787))))  severity failure;
	assert RAM(17788) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17788))))  severity failure;
	assert RAM(17789) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(17789))))  severity failure;
	assert RAM(17790) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17790))))  severity failure;
	assert RAM(17791) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17791))))  severity failure;
	assert RAM(17792) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(17792))))  severity failure;
	assert RAM(17793) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(17793))))  severity failure;
	assert RAM(17794) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17794))))  severity failure;
	assert RAM(17795) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17795))))  severity failure;
	assert RAM(17796) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17796))))  severity failure;
	assert RAM(17797) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17797))))  severity failure;
	assert RAM(17798) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17798))))  severity failure;
	assert RAM(17799) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17799))))  severity failure;
	assert RAM(17800) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17800))))  severity failure;
	assert RAM(17801) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(17801))))  severity failure;
	assert RAM(17802) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17802))))  severity failure;
	assert RAM(17803) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17803))))  severity failure;
	assert RAM(17804) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17804))))  severity failure;
	assert RAM(17805) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17805))))  severity failure;
	assert RAM(17806) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17806))))  severity failure;
	assert RAM(17807) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17807))))  severity failure;
	assert RAM(17808) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17808))))  severity failure;
	assert RAM(17809) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17809))))  severity failure;
	assert RAM(17810) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17810))))  severity failure;
	assert RAM(17811) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17811))))  severity failure;
	assert RAM(17812) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17812))))  severity failure;
	assert RAM(17813) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17813))))  severity failure;
	assert RAM(17814) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17814))))  severity failure;
	assert RAM(17815) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17815))))  severity failure;
	assert RAM(17816) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17816))))  severity failure;
	assert RAM(17817) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17817))))  severity failure;
	assert RAM(17818) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17818))))  severity failure;
	assert RAM(17819) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(17819))))  severity failure;
	assert RAM(17820) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17820))))  severity failure;
	assert RAM(17821) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17821))))  severity failure;
	assert RAM(17822) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17822))))  severity failure;
	assert RAM(17823) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17823))))  severity failure;
	assert RAM(17824) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17824))))  severity failure;
	assert RAM(17825) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17825))))  severity failure;
	assert RAM(17826) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17826))))  severity failure;
	assert RAM(17827) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(17827))))  severity failure;
	assert RAM(17828) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17828))))  severity failure;
	assert RAM(17829) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17829))))  severity failure;
	assert RAM(17830) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(17830))))  severity failure;
	assert RAM(17831) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17831))))  severity failure;
	assert RAM(17832) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17832))))  severity failure;
	assert RAM(17833) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17833))))  severity failure;
	assert RAM(17834) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17834))))  severity failure;
	assert RAM(17835) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17835))))  severity failure;
	assert RAM(17836) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17836))))  severity failure;
	assert RAM(17837) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17837))))  severity failure;
	assert RAM(17838) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17838))))  severity failure;
	assert RAM(17839) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17839))))  severity failure;
	assert RAM(17840) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17840))))  severity failure;
	assert RAM(17841) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17841))))  severity failure;
	assert RAM(17842) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17842))))  severity failure;
	assert RAM(17843) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17843))))  severity failure;
	assert RAM(17844) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17844))))  severity failure;
	assert RAM(17845) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17845))))  severity failure;
	assert RAM(17846) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17846))))  severity failure;
	assert RAM(17847) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17847))))  severity failure;
	assert RAM(17848) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17848))))  severity failure;
	assert RAM(17849) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(17849))))  severity failure;
	assert RAM(17850) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17850))))  severity failure;
	assert RAM(17851) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17851))))  severity failure;
	assert RAM(17852) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17852))))  severity failure;
	assert RAM(17853) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17853))))  severity failure;
	assert RAM(17854) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17854))))  severity failure;
	assert RAM(17855) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(17855))))  severity failure;
	assert RAM(17856) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17856))))  severity failure;
	assert RAM(17857) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17857))))  severity failure;
	assert RAM(17858) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17858))))  severity failure;
	assert RAM(17859) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17859))))  severity failure;
	assert RAM(17860) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17860))))  severity failure;
	assert RAM(17861) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17861))))  severity failure;
	assert RAM(17862) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17862))))  severity failure;
	assert RAM(17863) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17863))))  severity failure;
	assert RAM(17864) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(17864))))  severity failure;
	assert RAM(17865) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17865))))  severity failure;
	assert RAM(17866) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17866))))  severity failure;
	assert RAM(17867) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17867))))  severity failure;
	assert RAM(17868) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17868))))  severity failure;
	assert RAM(17869) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17869))))  severity failure;
	assert RAM(17870) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17870))))  severity failure;
	assert RAM(17871) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17871))))  severity failure;
	assert RAM(17872) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17872))))  severity failure;
	assert RAM(17873) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17873))))  severity failure;
	assert RAM(17874) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17874))))  severity failure;
	assert RAM(17875) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17875))))  severity failure;
	assert RAM(17876) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17876))))  severity failure;
	assert RAM(17877) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17877))))  severity failure;
	assert RAM(17878) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17878))))  severity failure;
	assert RAM(17879) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17879))))  severity failure;
	assert RAM(17880) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17880))))  severity failure;
	assert RAM(17881) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17881))))  severity failure;
	assert RAM(17882) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17882))))  severity failure;
	assert RAM(17883) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17883))))  severity failure;
	assert RAM(17884) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17884))))  severity failure;
	assert RAM(17885) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17885))))  severity failure;
	assert RAM(17886) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17886))))  severity failure;
	assert RAM(17887) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17887))))  severity failure;
	assert RAM(17888) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17888))))  severity failure;
	assert RAM(17889) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17889))))  severity failure;
	assert RAM(17890) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(17890))))  severity failure;
	assert RAM(17891) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17891))))  severity failure;
	assert RAM(17892) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17892))))  severity failure;
	assert RAM(17893) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17893))))  severity failure;
	assert RAM(17894) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17894))))  severity failure;
	assert RAM(17895) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17895))))  severity failure;
	assert RAM(17896) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17896))))  severity failure;
	assert RAM(17897) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(17897))))  severity failure;
	assert RAM(17898) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17898))))  severity failure;
	assert RAM(17899) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17899))))  severity failure;
	assert RAM(17900) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(17900))))  severity failure;
	assert RAM(17901) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17901))))  severity failure;
	assert RAM(17902) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17902))))  severity failure;
	assert RAM(17903) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17903))))  severity failure;
	assert RAM(17904) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17904))))  severity failure;
	assert RAM(17905) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17905))))  severity failure;
	assert RAM(17906) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17906))))  severity failure;
	assert RAM(17907) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17907))))  severity failure;
	assert RAM(17908) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(17908))))  severity failure;
	assert RAM(17909) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17909))))  severity failure;
	assert RAM(17910) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17910))))  severity failure;
	assert RAM(17911) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17911))))  severity failure;
	assert RAM(17912) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17912))))  severity failure;
	assert RAM(17913) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17913))))  severity failure;
	assert RAM(17914) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17914))))  severity failure;
	assert RAM(17915) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17915))))  severity failure;
	assert RAM(17916) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17916))))  severity failure;
	assert RAM(17917) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(17917))))  severity failure;
	assert RAM(17918) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17918))))  severity failure;
	assert RAM(17919) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17919))))  severity failure;
	assert RAM(17920) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17920))))  severity failure;
	assert RAM(17921) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17921))))  severity failure;
	assert RAM(17922) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(17922))))  severity failure;
	assert RAM(17923) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17923))))  severity failure;
	assert RAM(17924) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17924))))  severity failure;
	assert RAM(17925) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17925))))  severity failure;
	assert RAM(17926) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17926))))  severity failure;
	assert RAM(17927) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17927))))  severity failure;
	assert RAM(17928) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17928))))  severity failure;
	assert RAM(17929) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17929))))  severity failure;
	assert RAM(17930) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17930))))  severity failure;
	assert RAM(17931) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(17931))))  severity failure;
	assert RAM(17932) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17932))))  severity failure;
	assert RAM(17933) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(17933))))  severity failure;
	assert RAM(17934) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17934))))  severity failure;
	assert RAM(17935) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(17935))))  severity failure;
	assert RAM(17936) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17936))))  severity failure;
	assert RAM(17937) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17937))))  severity failure;
	assert RAM(17938) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17938))))  severity failure;
	assert RAM(17939) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17939))))  severity failure;
	assert RAM(17940) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17940))))  severity failure;
	assert RAM(17941) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17941))))  severity failure;
	assert RAM(17942) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17942))))  severity failure;
	assert RAM(17943) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17943))))  severity failure;
	assert RAM(17944) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17944))))  severity failure;
	assert RAM(17945) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17945))))  severity failure;
	assert RAM(17946) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(17946))))  severity failure;
	assert RAM(17947) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17947))))  severity failure;
	assert RAM(17948) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17948))))  severity failure;
	assert RAM(17949) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(17949))))  severity failure;
	assert RAM(17950) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(17950))))  severity failure;
	assert RAM(17951) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17951))))  severity failure;
	assert RAM(17952) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17952))))  severity failure;
	assert RAM(17953) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17953))))  severity failure;
	assert RAM(17954) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17954))))  severity failure;
	assert RAM(17955) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17955))))  severity failure;
	assert RAM(17956) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17956))))  severity failure;
	assert RAM(17957) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17957))))  severity failure;
	assert RAM(17958) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17958))))  severity failure;
	assert RAM(17959) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17959))))  severity failure;
	assert RAM(17960) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17960))))  severity failure;
	assert RAM(17961) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17961))))  severity failure;
	assert RAM(17962) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17962))))  severity failure;
	assert RAM(17963) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17963))))  severity failure;
	assert RAM(17964) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17964))))  severity failure;
	assert RAM(17965) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(17965))))  severity failure;
	assert RAM(17966) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17966))))  severity failure;
	assert RAM(17967) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17967))))  severity failure;
	assert RAM(17968) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17968))))  severity failure;
	assert RAM(17969) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17969))))  severity failure;
	assert RAM(17970) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17970))))  severity failure;
	assert RAM(17971) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17971))))  severity failure;
	assert RAM(17972) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17972))))  severity failure;
	assert RAM(17973) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(17973))))  severity failure;
	assert RAM(17974) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17974))))  severity failure;
	assert RAM(17975) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17975))))  severity failure;
	assert RAM(17976) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17976))))  severity failure;
	assert RAM(17977) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(17977))))  severity failure;
	assert RAM(17978) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(17978))))  severity failure;
	assert RAM(17979) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17979))))  severity failure;
	assert RAM(17980) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17980))))  severity failure;
	assert RAM(17981) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17981))))  severity failure;
	assert RAM(17982) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(17982))))  severity failure;
	assert RAM(17983) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17983))))  severity failure;
	assert RAM(17984) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17984))))  severity failure;
	assert RAM(17985) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17985))))  severity failure;
	assert RAM(17986) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17986))))  severity failure;
	assert RAM(17987) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17987))))  severity failure;
	assert RAM(17988) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17988))))  severity failure;
	assert RAM(17989) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17989))))  severity failure;
	assert RAM(17990) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17990))))  severity failure;
	assert RAM(17991) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17991))))  severity failure;
	assert RAM(17992) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17992))))  severity failure;
	assert RAM(17993) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17993))))  severity failure;
	assert RAM(17994) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17994))))  severity failure;
	assert RAM(17995) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17995))))  severity failure;
	assert RAM(17996) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17996))))  severity failure;
	assert RAM(17997) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17997))))  severity failure;
	assert RAM(17998) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17998))))  severity failure;
	assert RAM(17999) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17999))))  severity failure;
	assert RAM(18000) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18000))))  severity failure;
	assert RAM(18001) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18001))))  severity failure;
	assert RAM(18002) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18002))))  severity failure;
	assert RAM(18003) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18003))))  severity failure;
	assert RAM(18004) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18004))))  severity failure;
	assert RAM(18005) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18005))))  severity failure;
	assert RAM(18006) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18006))))  severity failure;
	assert RAM(18007) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18007))))  severity failure;
	assert RAM(18008) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(18008))))  severity failure;
	assert RAM(18009) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18009))))  severity failure;
	assert RAM(18010) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18010))))  severity failure;
	assert RAM(18011) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18011))))  severity failure;
	assert RAM(18012) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18012))))  severity failure;
	assert RAM(18013) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18013))))  severity failure;
	assert RAM(18014) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18014))))  severity failure;
	assert RAM(18015) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18015))))  severity failure;
	assert RAM(18016) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18016))))  severity failure;
	assert RAM(18017) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18017))))  severity failure;
	assert RAM(18018) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18018))))  severity failure;
	assert RAM(18019) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18019))))  severity failure;
	assert RAM(18020) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18020))))  severity failure;
	assert RAM(18021) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18021))))  severity failure;
	assert RAM(18022) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18022))))  severity failure;
	assert RAM(18023) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18023))))  severity failure;
	assert RAM(18024) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18024))))  severity failure;
	assert RAM(18025) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18025))))  severity failure;
	assert RAM(18026) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18026))))  severity failure;
	assert RAM(18027) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18027))))  severity failure;
	assert RAM(18028) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18028))))  severity failure;
	assert RAM(18029) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18029))))  severity failure;
	assert RAM(18030) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18030))))  severity failure;
	assert RAM(18031) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18031))))  severity failure;
	assert RAM(18032) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18032))))  severity failure;
	assert RAM(18033) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(18033))))  severity failure;
	assert RAM(18034) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18034))))  severity failure;
	assert RAM(18035) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18035))))  severity failure;
	assert RAM(18036) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(18036))))  severity failure;
	assert RAM(18037) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18037))))  severity failure;
	assert RAM(18038) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18038))))  severity failure;
	assert RAM(18039) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18039))))  severity failure;
	assert RAM(18040) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18040))))  severity failure;
	assert RAM(18041) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18041))))  severity failure;
	assert RAM(18042) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18042))))  severity failure;
	assert RAM(18043) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(18043))))  severity failure;
	assert RAM(18044) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18044))))  severity failure;
	assert RAM(18045) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18045))))  severity failure;
	assert RAM(18046) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18046))))  severity failure;
	assert RAM(18047) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18047))))  severity failure;
	assert RAM(18048) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18048))))  severity failure;
	assert RAM(18049) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18049))))  severity failure;
	assert RAM(18050) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(18050))))  severity failure;
	assert RAM(18051) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18051))))  severity failure;
	assert RAM(18052) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18052))))  severity failure;
	assert RAM(18053) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18053))))  severity failure;
	assert RAM(18054) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18054))))  severity failure;
	assert RAM(18055) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18055))))  severity failure;
	assert RAM(18056) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(18056))))  severity failure;
	assert RAM(18057) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18057))))  severity failure;
	assert RAM(18058) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18058))))  severity failure;
	assert RAM(18059) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18059))))  severity failure;
	assert RAM(18060) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18060))))  severity failure;
	assert RAM(18061) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18061))))  severity failure;
	assert RAM(18062) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18062))))  severity failure;
	assert RAM(18063) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18063))))  severity failure;
	assert RAM(18064) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18064))))  severity failure;
	assert RAM(18065) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(18065))))  severity failure;
	assert RAM(18066) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18066))))  severity failure;
	assert RAM(18067) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18067))))  severity failure;
	assert RAM(18068) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18068))))  severity failure;
	assert RAM(18069) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18069))))  severity failure;
	assert RAM(18070) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18070))))  severity failure;
	assert RAM(18071) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(18071))))  severity failure;
	assert RAM(18072) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18072))))  severity failure;
	assert RAM(18073) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18073))))  severity failure;
	assert RAM(18074) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18074))))  severity failure;
	assert RAM(18075) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18075))))  severity failure;
	assert RAM(18076) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18076))))  severity failure;
	assert RAM(18077) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18077))))  severity failure;
	assert RAM(18078) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18078))))  severity failure;
	assert RAM(18079) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18079))))  severity failure;
	assert RAM(18080) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18080))))  severity failure;
	assert RAM(18081) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18081))))  severity failure;
	assert RAM(18082) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18082))))  severity failure;
	assert RAM(18083) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18083))))  severity failure;
	assert RAM(18084) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18084))))  severity failure;
	assert RAM(18085) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18085))))  severity failure;
	assert RAM(18086) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18086))))  severity failure;
	assert RAM(18087) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18087))))  severity failure;
	assert RAM(18088) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(18088))))  severity failure;
	assert RAM(18089) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18089))))  severity failure;
	assert RAM(18090) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18090))))  severity failure;
	assert RAM(18091) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18091))))  severity failure;
	assert RAM(18092) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18092))))  severity failure;
	assert RAM(18093) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18093))))  severity failure;
	assert RAM(18094) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18094))))  severity failure;
	assert RAM(18095) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18095))))  severity failure;
	assert RAM(18096) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18096))))  severity failure;
	assert RAM(18097) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18097))))  severity failure;
	assert RAM(18098) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18098))))  severity failure;
	assert RAM(18099) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18099))))  severity failure;
	assert RAM(18100) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(18100))))  severity failure;
	assert RAM(18101) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18101))))  severity failure;
	assert RAM(18102) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18102))))  severity failure;
	assert RAM(18103) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18103))))  severity failure;
	assert RAM(18104) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18104))))  severity failure;
	assert RAM(18105) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18105))))  severity failure;
	assert RAM(18106) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18106))))  severity failure;
	assert RAM(18107) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(18107))))  severity failure;
	assert RAM(18108) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18108))))  severity failure;
	assert RAM(18109) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18109))))  severity failure;
	assert RAM(18110) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18110))))  severity failure;
	assert RAM(18111) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18111))))  severity failure;
	assert RAM(18112) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18112))))  severity failure;
	assert RAM(18113) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18113))))  severity failure;
	assert RAM(18114) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18114))))  severity failure;
	assert RAM(18115) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18115))))  severity failure;
	assert RAM(18116) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18116))))  severity failure;
	assert RAM(18117) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18117))))  severity failure;
	assert RAM(18118) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18118))))  severity failure;
	assert RAM(18119) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(18119))))  severity failure;
	assert RAM(18120) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(18120))))  severity failure;
	assert RAM(18121) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(18121))))  severity failure;
	assert RAM(18122) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18122))))  severity failure;
	assert RAM(18123) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18123))))  severity failure;
	assert RAM(18124) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(18124))))  severity failure;
	assert RAM(18125) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18125))))  severity failure;
	assert RAM(18126) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18126))))  severity failure;
	assert RAM(18127) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18127))))  severity failure;
	assert RAM(18128) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18128))))  severity failure;
	assert RAM(18129) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18129))))  severity failure;
	assert RAM(18130) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18130))))  severity failure;
	assert RAM(18131) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18131))))  severity failure;
	assert RAM(18132) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18132))))  severity failure;
	assert RAM(18133) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18133))))  severity failure;
	assert RAM(18134) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18134))))  severity failure;
	assert RAM(18135) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(18135))))  severity failure;
	assert RAM(18136) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(18136))))  severity failure;
	assert RAM(18137) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18137))))  severity failure;
	assert RAM(18138) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(18138))))  severity failure;
	assert RAM(18139) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18139))))  severity failure;
	assert RAM(18140) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18140))))  severity failure;
	assert RAM(18141) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18141))))  severity failure;
	assert RAM(18142) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18142))))  severity failure;
	assert RAM(18143) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(18143))))  severity failure;
	assert RAM(18144) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18144))))  severity failure;
	assert RAM(18145) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18145))))  severity failure;
	assert RAM(18146) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18146))))  severity failure;
	assert RAM(18147) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18147))))  severity failure;
	assert RAM(18148) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18148))))  severity failure;
	assert RAM(18149) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18149))))  severity failure;
	assert RAM(18150) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18150))))  severity failure;
	assert RAM(18151) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(18151))))  severity failure;
	assert RAM(18152) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18152))))  severity failure;
	assert RAM(18153) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18153))))  severity failure;
	assert RAM(18154) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18154))))  severity failure;
	assert RAM(18155) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18155))))  severity failure;
	assert RAM(18156) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18156))))  severity failure;
	assert RAM(18157) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18157))))  severity failure;
	assert RAM(18158) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18158))))  severity failure;
	assert RAM(18159) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(18159))))  severity failure;
	assert RAM(18160) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18160))))  severity failure;
	assert RAM(18161) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18161))))  severity failure;
	assert RAM(18162) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18162))))  severity failure;
	assert RAM(18163) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18163))))  severity failure;
	assert RAM(18164) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18164))))  severity failure;
	assert RAM(18165) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18165))))  severity failure;
	assert RAM(18166) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18166))))  severity failure;
	assert RAM(18167) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18167))))  severity failure;
	assert RAM(18168) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18168))))  severity failure;
	assert RAM(18169) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18169))))  severity failure;
	assert RAM(18170) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18170))))  severity failure;
	assert RAM(18171) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18171))))  severity failure;
	assert RAM(18172) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18172))))  severity failure;
	assert RAM(18173) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18173))))  severity failure;
	assert RAM(18174) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18174))))  severity failure;
	assert RAM(18175) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18175))))  severity failure;
	assert RAM(18176) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18176))))  severity failure;
	assert RAM(18177) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18177))))  severity failure;
	assert RAM(18178) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18178))))  severity failure;
	assert RAM(18179) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18179))))  severity failure;
	assert RAM(18180) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(18180))))  severity failure;
	assert RAM(18181) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18181))))  severity failure;
	assert RAM(18182) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18182))))  severity failure;
	assert RAM(18183) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18183))))  severity failure;
	assert RAM(18184) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18184))))  severity failure;
	assert RAM(18185) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18185))))  severity failure;
	assert RAM(18186) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18186))))  severity failure;
	assert RAM(18187) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18187))))  severity failure;
	assert RAM(18188) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18188))))  severity failure;
	assert RAM(18189) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18189))))  severity failure;
	assert RAM(18190) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18190))))  severity failure;
	assert RAM(18191) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18191))))  severity failure;
	assert RAM(18192) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18192))))  severity failure;
	assert RAM(18193) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18193))))  severity failure;
	assert RAM(18194) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18194))))  severity failure;
	assert RAM(18195) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18195))))  severity failure;
	assert RAM(18196) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18196))))  severity failure;
	assert RAM(18197) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18197))))  severity failure;
	assert RAM(18198) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18198))))  severity failure;
	assert RAM(18199) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18199))))  severity failure;
	assert RAM(18200) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18200))))  severity failure;
	assert RAM(18201) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18201))))  severity failure;
	assert RAM(18202) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18202))))  severity failure;
	assert RAM(18203) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(18203))))  severity failure;
	assert RAM(18204) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18204))))  severity failure;
	assert RAM(18205) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18205))))  severity failure;
	assert RAM(18206) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(18206))))  severity failure;
	assert RAM(18207) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18207))))  severity failure;
	assert RAM(18208) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(18208))))  severity failure;
	assert RAM(18209) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18209))))  severity failure;
	assert RAM(18210) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(18210))))  severity failure;
	assert RAM(18211) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18211))))  severity failure;
	assert RAM(18212) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18212))))  severity failure;
	assert RAM(18213) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18213))))  severity failure;
	assert RAM(18214) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18214))))  severity failure;
	assert RAM(18215) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18215))))  severity failure;
	assert RAM(18216) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18216))))  severity failure;
	assert RAM(18217) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18217))))  severity failure;
	assert RAM(18218) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(18218))))  severity failure;
	assert RAM(18219) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18219))))  severity failure;
	assert RAM(18220) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18220))))  severity failure;
	assert RAM(18221) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18221))))  severity failure;
	assert RAM(18222) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18222))))  severity failure;
	assert RAM(18223) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18223))))  severity failure;
	assert RAM(18224) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18224))))  severity failure;
	assert RAM(18225) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18225))))  severity failure;
	assert RAM(18226) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18226))))  severity failure;
	assert RAM(18227) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18227))))  severity failure;
	assert RAM(18228) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18228))))  severity failure;
	assert RAM(18229) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18229))))  severity failure;
	assert RAM(18230) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18230))))  severity failure;
	assert RAM(18231) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18231))))  severity failure;
	assert RAM(18232) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(18232))))  severity failure;
	assert RAM(18233) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18233))))  severity failure;
	assert RAM(18234) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18234))))  severity failure;
	assert RAM(18235) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(18235))))  severity failure;
	assert RAM(18236) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18236))))  severity failure;
	assert RAM(18237) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18237))))  severity failure;
	assert RAM(18238) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18238))))  severity failure;
	assert RAM(18239) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18239))))  severity failure;
	assert RAM(18240) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(18240))))  severity failure;
	assert RAM(18241) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18241))))  severity failure;
	assert RAM(18242) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18242))))  severity failure;
	assert RAM(18243) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18243))))  severity failure;
	assert RAM(18244) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18244))))  severity failure;
	assert RAM(18245) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18245))))  severity failure;
	assert RAM(18246) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18246))))  severity failure;
	assert RAM(18247) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18247))))  severity failure;
	assert RAM(18248) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(18248))))  severity failure;
	assert RAM(18249) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18249))))  severity failure;
	assert RAM(18250) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18250))))  severity failure;
	assert RAM(18251) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18251))))  severity failure;
	assert RAM(18252) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18252))))  severity failure;
	assert RAM(18253) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18253))))  severity failure;
	assert RAM(18254) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18254))))  severity failure;
	assert RAM(18255) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(18255))))  severity failure;
	assert RAM(18256) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(18256))))  severity failure;
	assert RAM(18257) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18257))))  severity failure;
	assert RAM(18258) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18258))))  severity failure;
	assert RAM(18259) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18259))))  severity failure;
	assert RAM(18260) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18260))))  severity failure;
	assert RAM(18261) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18261))))  severity failure;
	assert RAM(18262) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18262))))  severity failure;
	assert RAM(18263) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18263))))  severity failure;
	assert RAM(18264) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18264))))  severity failure;
	assert RAM(18265) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18265))))  severity failure;
	assert RAM(18266) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18266))))  severity failure;
	assert RAM(18267) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18267))))  severity failure;
	assert RAM(18268) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18268))))  severity failure;
	assert RAM(18269) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18269))))  severity failure;
	assert RAM(18270) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18270))))  severity failure;
	assert RAM(18271) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(18271))))  severity failure;
	assert RAM(18272) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18272))))  severity failure;
	assert RAM(18273) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18273))))  severity failure;
	assert RAM(18274) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18274))))  severity failure;
	assert RAM(18275) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18275))))  severity failure;
	assert RAM(18276) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18276))))  severity failure;
	assert RAM(18277) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18277))))  severity failure;
	assert RAM(18278) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18278))))  severity failure;
	assert RAM(18279) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18279))))  severity failure;
	assert RAM(18280) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(18280))))  severity failure;
	assert RAM(18281) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18281))))  severity failure;
	assert RAM(18282) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(18282))))  severity failure;
	assert RAM(18283) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18283))))  severity failure;
	assert RAM(18284) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18284))))  severity failure;
	assert RAM(18285) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(18285))))  severity failure;
	assert RAM(18286) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(18286))))  severity failure;
	assert RAM(18287) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18287))))  severity failure;
	assert RAM(18288) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18288))))  severity failure;
	assert RAM(18289) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18289))))  severity failure;
	assert RAM(18290) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18290))))  severity failure;
	assert RAM(18291) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18291))))  severity failure;
	assert RAM(18292) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18292))))  severity failure;
	assert RAM(18293) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18293))))  severity failure;
	assert RAM(18294) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18294))))  severity failure;
	assert RAM(18295) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18295))))  severity failure;
	assert RAM(18296) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18296))))  severity failure;
	assert RAM(18297) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18297))))  severity failure;
	assert RAM(18298) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(18298))))  severity failure;
	assert RAM(18299) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18299))))  severity failure;
	assert RAM(18300) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18300))))  severity failure;
	assert RAM(18301) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18301))))  severity failure;
	assert RAM(18302) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18302))))  severity failure;
	assert RAM(18303) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18303))))  severity failure;
	assert RAM(18304) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18304))))  severity failure;
	assert RAM(18305) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18305))))  severity failure;
	assert RAM(18306) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18306))))  severity failure;
	assert RAM(18307) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18307))))  severity failure;
	assert RAM(18308) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18308))))  severity failure;
	assert RAM(18309) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18309))))  severity failure;
	assert RAM(18310) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18310))))  severity failure;
	assert RAM(18311) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18311))))  severity failure;
	assert RAM(18312) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(18312))))  severity failure;
	assert RAM(18313) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18313))))  severity failure;
	assert RAM(18314) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18314))))  severity failure;
	assert RAM(18315) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18315))))  severity failure;
	assert RAM(18316) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18316))))  severity failure;
	assert RAM(18317) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18317))))  severity failure;
	assert RAM(18318) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18318))))  severity failure;
	assert RAM(18319) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18319))))  severity failure;
	assert RAM(18320) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18320))))  severity failure;
	assert RAM(18321) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18321))))  severity failure;
	assert RAM(18322) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18322))))  severity failure;
	assert RAM(18323) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18323))))  severity failure;
	assert RAM(18324) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18324))))  severity failure;
	assert RAM(18325) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(18325))))  severity failure;
	assert RAM(18326) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18326))))  severity failure;
	assert RAM(18327) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18327))))  severity failure;
	assert RAM(18328) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18328))))  severity failure;
	assert RAM(18329) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18329))))  severity failure;
	assert RAM(18330) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18330))))  severity failure;
	assert RAM(18331) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18331))))  severity failure;
	assert RAM(18332) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18332))))  severity failure;
	assert RAM(18333) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18333))))  severity failure;
	assert RAM(18334) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18334))))  severity failure;
	assert RAM(18335) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18335))))  severity failure;
	assert RAM(18336) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18336))))  severity failure;
	assert RAM(18337) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18337))))  severity failure;
	assert RAM(18338) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(18338))))  severity failure;
	assert RAM(18339) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18339))))  severity failure;
	assert RAM(18340) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(18340))))  severity failure;
	assert RAM(18341) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18341))))  severity failure;
	assert RAM(18342) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18342))))  severity failure;
	assert RAM(18343) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18343))))  severity failure;
	assert RAM(18344) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(18344))))  severity failure;
	assert RAM(18345) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18345))))  severity failure;
	assert RAM(18346) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18346))))  severity failure;
	assert RAM(18347) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18347))))  severity failure;
	assert RAM(18348) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18348))))  severity failure;
	assert RAM(18349) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18349))))  severity failure;
	assert RAM(18350) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18350))))  severity failure;
	assert RAM(18351) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18351))))  severity failure;
	assert RAM(18352) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18352))))  severity failure;
	assert RAM(18353) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18353))))  severity failure;
	assert RAM(18354) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18354))))  severity failure;
	assert RAM(18355) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18355))))  severity failure;
	assert RAM(18356) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18356))))  severity failure;
	assert RAM(18357) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18357))))  severity failure;
	assert RAM(18358) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(18358))))  severity failure;
	assert RAM(18359) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18359))))  severity failure;
	assert RAM(18360) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18360))))  severity failure;
	assert RAM(18361) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18361))))  severity failure;
	assert RAM(18362) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18362))))  severity failure;
	assert RAM(18363) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18363))))  severity failure;
	assert RAM(18364) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18364))))  severity failure;
	assert RAM(18365) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18365))))  severity failure;
	assert RAM(18366) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18366))))  severity failure;
	assert RAM(18367) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18367))))  severity failure;
	assert RAM(18368) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18368))))  severity failure;
	assert RAM(18369) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18369))))  severity failure;
	assert RAM(18370) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18370))))  severity failure;
	assert RAM(18371) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18371))))  severity failure;
	assert RAM(18372) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18372))))  severity failure;
	assert RAM(18373) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18373))))  severity failure;
	assert RAM(18374) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18374))))  severity failure;
	assert RAM(18375) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18375))))  severity failure;
	assert RAM(18376) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18376))))  severity failure;
	assert RAM(18377) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18377))))  severity failure;
	assert RAM(18378) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18378))))  severity failure;
	assert RAM(18379) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18379))))  severity failure;
	assert RAM(18380) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18380))))  severity failure;
	assert RAM(18381) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18381))))  severity failure;
	assert RAM(18382) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18382))))  severity failure;
	assert RAM(18383) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18383))))  severity failure;
	assert RAM(18384) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18384))))  severity failure;
	assert RAM(18385) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18385))))  severity failure;
	assert RAM(18386) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18386))))  severity failure;
	assert RAM(18387) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18387))))  severity failure;
	assert RAM(18388) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18388))))  severity failure;
	assert RAM(18389) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18389))))  severity failure;
	assert RAM(18390) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18390))))  severity failure;
	assert RAM(18391) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(18391))))  severity failure;
	assert RAM(18392) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18392))))  severity failure;
	assert RAM(18393) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18393))))  severity failure;
	assert RAM(18394) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18394))))  severity failure;
	assert RAM(18395) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18395))))  severity failure;
	assert RAM(18396) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18396))))  severity failure;
	assert RAM(18397) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(18397))))  severity failure;
	assert RAM(18398) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18398))))  severity failure;
	assert RAM(18399) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18399))))  severity failure;
	assert RAM(18400) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18400))))  severity failure;
	assert RAM(18401) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18401))))  severity failure;
	assert RAM(18402) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18402))))  severity failure;
	assert RAM(18403) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18403))))  severity failure;
	assert RAM(18404) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(18404))))  severity failure;
	assert RAM(18405) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18405))))  severity failure;
	assert RAM(18406) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18406))))  severity failure;
	assert RAM(18407) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(18407))))  severity failure;
	assert RAM(18408) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18408))))  severity failure;
	assert RAM(18409) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18409))))  severity failure;
	assert RAM(18410) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(18410))))  severity failure;
	assert RAM(18411) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18411))))  severity failure;
	assert RAM(18412) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18412))))  severity failure;
	assert RAM(18413) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18413))))  severity failure;
	assert RAM(18414) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18414))))  severity failure;
	assert RAM(18415) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18415))))  severity failure;
	assert RAM(18416) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18416))))  severity failure;
	assert RAM(18417) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18417))))  severity failure;
	assert RAM(18418) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18418))))  severity failure;
	assert RAM(18419) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18419))))  severity failure;
	assert RAM(18420) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18420))))  severity failure;
	assert RAM(18421) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18421))))  severity failure;
	assert RAM(18422) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18422))))  severity failure;
	assert RAM(18423) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18423))))  severity failure;
	assert RAM(18424) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(18424))))  severity failure;
	assert RAM(18425) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18425))))  severity failure;
	assert RAM(18426) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18426))))  severity failure;
	assert RAM(18427) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18427))))  severity failure;
	assert RAM(18428) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18428))))  severity failure;
	assert RAM(18429) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18429))))  severity failure;
	assert RAM(18430) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18430))))  severity failure;
	assert RAM(18431) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18431))))  severity failure;
	assert RAM(18432) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(18432))))  severity failure;
	assert RAM(18433) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(18433))))  severity failure;
	assert RAM(18434) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18434))))  severity failure;
	assert RAM(18435) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18435))))  severity failure;
	assert RAM(18436) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18436))))  severity failure;
	assert RAM(18437) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18437))))  severity failure;
	assert RAM(18438) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18438))))  severity failure;
	assert RAM(18439) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18439))))  severity failure;
	assert RAM(18440) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18440))))  severity failure;
	assert RAM(18441) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18441))))  severity failure;
	assert RAM(18442) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(18442))))  severity failure;
	assert RAM(18443) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18443))))  severity failure;
	assert RAM(18444) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18444))))  severity failure;
	assert RAM(18445) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(18445))))  severity failure;
	assert RAM(18446) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18446))))  severity failure;
	assert RAM(18447) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18447))))  severity failure;
	assert RAM(18448) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18448))))  severity failure;
	assert RAM(18449) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18449))))  severity failure;
	assert RAM(18450) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18450))))  severity failure;
	assert RAM(18451) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18451))))  severity failure;
	assert RAM(18452) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18452))))  severity failure;
	assert RAM(18453) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18453))))  severity failure;
	assert RAM(18454) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18454))))  severity failure;
	assert RAM(18455) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18455))))  severity failure;
	assert RAM(18456) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18456))))  severity failure;
	assert RAM(18457) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(18457))))  severity failure;
	assert RAM(18458) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18458))))  severity failure;
	assert RAM(18459) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18459))))  severity failure;
	assert RAM(18460) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18460))))  severity failure;
	assert RAM(18461) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18461))))  severity failure;
	assert RAM(18462) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18462))))  severity failure;
	assert RAM(18463) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18463))))  severity failure;
	assert RAM(18464) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18464))))  severity failure;
	assert RAM(18465) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18465))))  severity failure;
	assert RAM(18466) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18466))))  severity failure;
	assert RAM(18467) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18467))))  severity failure;
	assert RAM(18468) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18468))))  severity failure;
	assert RAM(18469) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18469))))  severity failure;
	assert RAM(18470) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18470))))  severity failure;
	assert RAM(18471) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18471))))  severity failure;
	assert RAM(18472) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18472))))  severity failure;
	assert RAM(18473) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18473))))  severity failure;
	assert RAM(18474) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18474))))  severity failure;
	assert RAM(18475) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18475))))  severity failure;
	assert RAM(18476) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18476))))  severity failure;
	assert RAM(18477) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(18477))))  severity failure;
	assert RAM(18478) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18478))))  severity failure;
	assert RAM(18479) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(18479))))  severity failure;
	assert RAM(18480) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18480))))  severity failure;
	assert RAM(18481) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18481))))  severity failure;
	assert RAM(18482) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18482))))  severity failure;
	assert RAM(18483) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18483))))  severity failure;
	assert RAM(18484) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18484))))  severity failure;
	assert RAM(18485) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18485))))  severity failure;
	assert RAM(18486) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18486))))  severity failure;
	assert RAM(18487) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18487))))  severity failure;
	assert RAM(18488) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18488))))  severity failure;
	assert RAM(18489) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(18489))))  severity failure;
	assert RAM(18490) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18490))))  severity failure;
	assert RAM(18491) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18491))))  severity failure;
	assert RAM(18492) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18492))))  severity failure;
	assert RAM(18493) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(18493))))  severity failure;
	assert RAM(18494) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18494))))  severity failure;
	assert RAM(18495) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18495))))  severity failure;
	assert RAM(18496) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18496))))  severity failure;
	assert RAM(18497) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18497))))  severity failure;
	assert RAM(18498) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18498))))  severity failure;
	assert RAM(18499) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18499))))  severity failure;
	assert RAM(18500) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18500))))  severity failure;
	assert RAM(18501) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18501))))  severity failure;
	assert RAM(18502) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18502))))  severity failure;
	assert RAM(18503) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(18503))))  severity failure;
	assert RAM(18504) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18504))))  severity failure;
	assert RAM(18505) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18505))))  severity failure;
	assert RAM(18506) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18506))))  severity failure;
	assert RAM(18507) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18507))))  severity failure;
	assert RAM(18508) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18508))))  severity failure;
	assert RAM(18509) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18509))))  severity failure;
	assert RAM(18510) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18510))))  severity failure;
	assert RAM(18511) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(18511))))  severity failure;
	assert RAM(18512) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18512))))  severity failure;
	assert RAM(18513) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18513))))  severity failure;
	assert RAM(18514) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(18514))))  severity failure;
	assert RAM(18515) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18515))))  severity failure;
	assert RAM(18516) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18516))))  severity failure;
	assert RAM(18517) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18517))))  severity failure;
	assert RAM(18518) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18518))))  severity failure;
	assert RAM(18519) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18519))))  severity failure;
	assert RAM(18520) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18520))))  severity failure;
	assert RAM(18521) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18521))))  severity failure;
	assert RAM(18522) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18522))))  severity failure;
	assert RAM(18523) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18523))))  severity failure;
	assert RAM(18524) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18524))))  severity failure;
	assert RAM(18525) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18525))))  severity failure;
	assert RAM(18526) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18526))))  severity failure;
	assert RAM(18527) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18527))))  severity failure;
	assert RAM(18528) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18528))))  severity failure;
	assert RAM(18529) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18529))))  severity failure;
	assert RAM(18530) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18530))))  severity failure;
	assert RAM(18531) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(18531))))  severity failure;
	assert RAM(18532) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18532))))  severity failure;
	assert RAM(18533) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18533))))  severity failure;
	assert RAM(18534) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18534))))  severity failure;
	assert RAM(18535) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(18535))))  severity failure;
	assert RAM(18536) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18536))))  severity failure;
	assert RAM(18537) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18537))))  severity failure;
	assert RAM(18538) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18538))))  severity failure;
	assert RAM(18539) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18539))))  severity failure;
	assert RAM(18540) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18540))))  severity failure;
	assert RAM(18541) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18541))))  severity failure;
	assert RAM(18542) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18542))))  severity failure;
	assert RAM(18543) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18543))))  severity failure;
	assert RAM(18544) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(18544))))  severity failure;
	assert RAM(18545) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18545))))  severity failure;
	assert RAM(18546) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18546))))  severity failure;
	assert RAM(18547) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18547))))  severity failure;
	assert RAM(18548) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18548))))  severity failure;
	assert RAM(18549) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18549))))  severity failure;
	assert RAM(18550) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18550))))  severity failure;
	assert RAM(18551) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18551))))  severity failure;
	assert RAM(18552) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18552))))  severity failure;
	assert RAM(18553) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18553))))  severity failure;
	assert RAM(18554) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18554))))  severity failure;
	assert RAM(18555) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18555))))  severity failure;
	assert RAM(18556) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18556))))  severity failure;
	assert RAM(18557) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18557))))  severity failure;
	assert RAM(18558) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18558))))  severity failure;
	assert RAM(18559) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18559))))  severity failure;
	assert RAM(18560) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18560))))  severity failure;
	assert RAM(18561) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18561))))  severity failure;
	assert RAM(18562) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18562))))  severity failure;
	assert RAM(18563) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18563))))  severity failure;
	assert RAM(18564) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18564))))  severity failure;
	assert RAM(18565) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18565))))  severity failure;
	assert RAM(18566) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18566))))  severity failure;
	assert RAM(18567) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18567))))  severity failure;
	assert RAM(18568) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18568))))  severity failure;
	assert RAM(18569) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18569))))  severity failure;
	assert RAM(18570) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18570))))  severity failure;
	assert RAM(18571) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18571))))  severity failure;
	assert RAM(18572) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18572))))  severity failure;
	assert RAM(18573) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18573))))  severity failure;
	assert RAM(18574) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18574))))  severity failure;
	assert RAM(18575) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18575))))  severity failure;
	assert RAM(18576) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(18576))))  severity failure;
	assert RAM(18577) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18577))))  severity failure;
	assert RAM(18578) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18578))))  severity failure;
	assert RAM(18579) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18579))))  severity failure;
	assert RAM(18580) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18580))))  severity failure;
	assert RAM(18581) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18581))))  severity failure;
	assert RAM(18582) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18582))))  severity failure;
	assert RAM(18583) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18583))))  severity failure;
	assert RAM(18584) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18584))))  severity failure;
	assert RAM(18585) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18585))))  severity failure;
	assert RAM(18586) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18586))))  severity failure;
	assert RAM(18587) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18587))))  severity failure;
	assert RAM(18588) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(18588))))  severity failure;
	assert RAM(18589) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18589))))  severity failure;
	assert RAM(18590) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18590))))  severity failure;
	assert RAM(18591) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18591))))  severity failure;
	assert RAM(18592) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18592))))  severity failure;
	assert RAM(18593) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(18593))))  severity failure;
	assert RAM(18594) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18594))))  severity failure;
	assert RAM(18595) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18595))))  severity failure;
	assert RAM(18596) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18596))))  severity failure;
	assert RAM(18597) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(18597))))  severity failure;
	assert RAM(18598) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18598))))  severity failure;
	assert RAM(18599) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18599))))  severity failure;
	assert RAM(18600) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18600))))  severity failure;
	assert RAM(18601) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18601))))  severity failure;
	assert RAM(18602) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18602))))  severity failure;
	assert RAM(18603) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18603))))  severity failure;
	assert RAM(18604) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18604))))  severity failure;
	assert RAM(18605) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18605))))  severity failure;
	assert RAM(18606) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18606))))  severity failure;
	assert RAM(18607) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18607))))  severity failure;
	assert RAM(18608) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18608))))  severity failure;
	assert RAM(18609) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18609))))  severity failure;
	assert RAM(18610) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18610))))  severity failure;
	assert RAM(18611) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18611))))  severity failure;
	assert RAM(18612) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18612))))  severity failure;
	assert RAM(18613) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18613))))  severity failure;
	assert RAM(18614) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(18614))))  severity failure;
	assert RAM(18615) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18615))))  severity failure;
	assert RAM(18616) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18616))))  severity failure;
	assert RAM(18617) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18617))))  severity failure;
	assert RAM(18618) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18618))))  severity failure;
	assert RAM(18619) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18619))))  severity failure;
	assert RAM(18620) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18620))))  severity failure;
	assert RAM(18621) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18621))))  severity failure;
	assert RAM(18622) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(18622))))  severity failure;
	assert RAM(18623) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18623))))  severity failure;
	assert RAM(18624) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(18624))))  severity failure;
	assert RAM(18625) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18625))))  severity failure;
	assert RAM(18626) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18626))))  severity failure;
	assert RAM(18627) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18627))))  severity failure;
	assert RAM(18628) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18628))))  severity failure;
	assert RAM(18629) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18629))))  severity failure;
	assert RAM(18630) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18630))))  severity failure;
	assert RAM(18631) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18631))))  severity failure;
	assert RAM(18632) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18632))))  severity failure;
	assert RAM(18633) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18633))))  severity failure;
	assert RAM(18634) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18634))))  severity failure;
	assert RAM(18635) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18635))))  severity failure;
	assert RAM(18636) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18636))))  severity failure;
	assert RAM(18637) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18637))))  severity failure;
	assert RAM(18638) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18638))))  severity failure;
	assert RAM(18639) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18639))))  severity failure;
	assert RAM(18640) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18640))))  severity failure;
	assert RAM(18641) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18641))))  severity failure;
	assert RAM(18642) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18642))))  severity failure;
	assert RAM(18643) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18643))))  severity failure;
	assert RAM(18644) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18644))))  severity failure;
	assert RAM(18645) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18645))))  severity failure;
	assert RAM(18646) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18646))))  severity failure;
	assert RAM(18647) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18647))))  severity failure;
	assert RAM(18648) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(18648))))  severity failure;
	assert RAM(18649) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18649))))  severity failure;
	assert RAM(18650) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18650))))  severity failure;
	assert RAM(18651) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18651))))  severity failure;
	assert RAM(18652) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(18652))))  severity failure;
	assert RAM(18653) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(18653))))  severity failure;
	assert RAM(18654) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18654))))  severity failure;
	assert RAM(18655) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18655))))  severity failure;
	assert RAM(18656) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18656))))  severity failure;
	assert RAM(18657) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18657))))  severity failure;
	assert RAM(18658) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18658))))  severity failure;
	assert RAM(18659) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18659))))  severity failure;
	assert RAM(18660) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(18660))))  severity failure;
	assert RAM(18661) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(18661))))  severity failure;
	assert RAM(18662) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(18662))))  severity failure;
	assert RAM(18663) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18663))))  severity failure;
	assert RAM(18664) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18664))))  severity failure;
	assert RAM(18665) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18665))))  severity failure;
	assert RAM(18666) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(18666))))  severity failure;
	assert RAM(18667) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18667))))  severity failure;
	assert RAM(18668) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(18668))))  severity failure;
	assert RAM(18669) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18669))))  severity failure;
	assert RAM(18670) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18670))))  severity failure;
	assert RAM(18671) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18671))))  severity failure;
	assert RAM(18672) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18672))))  severity failure;
	assert RAM(18673) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18673))))  severity failure;
	assert RAM(18674) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18674))))  severity failure;
	assert RAM(18675) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18675))))  severity failure;
	assert RAM(18676) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(18676))))  severity failure;
	assert RAM(18677) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18677))))  severity failure;
	assert RAM(18678) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18678))))  severity failure;
	assert RAM(18679) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18679))))  severity failure;
	assert RAM(18680) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(18680))))  severity failure;
	assert RAM(18681) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18681))))  severity failure;
	assert RAM(18682) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18682))))  severity failure;
	assert RAM(18683) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18683))))  severity failure;
	assert RAM(18684) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18684))))  severity failure;
	assert RAM(18685) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18685))))  severity failure;
	assert RAM(18686) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18686))))  severity failure;
	assert RAM(18687) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18687))))  severity failure;
	assert RAM(18688) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18688))))  severity failure;
	assert RAM(18689) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18689))))  severity failure;
	assert RAM(18690) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18690))))  severity failure;
	assert RAM(18691) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18691))))  severity failure;
	assert RAM(18692) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18692))))  severity failure;
	assert RAM(18693) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18693))))  severity failure;
	assert RAM(18694) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18694))))  severity failure;
	assert RAM(18695) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18695))))  severity failure;
	assert RAM(18696) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18696))))  severity failure;
	assert RAM(18697) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18697))))  severity failure;
	assert RAM(18698) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18698))))  severity failure;
	assert RAM(18699) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18699))))  severity failure;
	assert RAM(18700) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18700))))  severity failure;
	assert RAM(18701) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18701))))  severity failure;
	assert RAM(18702) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(18702))))  severity failure;
	assert RAM(18703) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18703))))  severity failure;
	assert RAM(18704) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18704))))  severity failure;
	assert RAM(18705) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(18705))))  severity failure;
	assert RAM(18706) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18706))))  severity failure;
	assert RAM(18707) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(18707))))  severity failure;
	assert RAM(18708) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18708))))  severity failure;
	assert RAM(18709) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18709))))  severity failure;
	assert RAM(18710) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(18710))))  severity failure;
	assert RAM(18711) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18711))))  severity failure;
	assert RAM(18712) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(18712))))  severity failure;
	assert RAM(18713) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(18713))))  severity failure;
	assert RAM(18714) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18714))))  severity failure;
	assert RAM(18715) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(18715))))  severity failure;
	assert RAM(18716) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(18716))))  severity failure;
	assert RAM(18717) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18717))))  severity failure;
	assert RAM(18718) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(18718))))  severity failure;
	assert RAM(18719) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18719))))  severity failure;
	assert RAM(18720) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18720))))  severity failure;
	assert RAM(18721) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(18721))))  severity failure;
	assert RAM(18722) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18722))))  severity failure;
	assert RAM(18723) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18723))))  severity failure;
	assert RAM(18724) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18724))))  severity failure;
	assert RAM(18725) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18725))))  severity failure;
	assert RAM(18726) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18726))))  severity failure;
	assert RAM(18727) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18727))))  severity failure;
	assert RAM(18728) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18728))))  severity failure;
	assert RAM(18729) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18729))))  severity failure;
	assert RAM(18730) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18730))))  severity failure;
	assert RAM(18731) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18731))))  severity failure;
	assert RAM(18732) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18732))))  severity failure;
	assert RAM(18733) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18733))))  severity failure;
	assert RAM(18734) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18734))))  severity failure;
	assert RAM(18735) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18735))))  severity failure;
	assert RAM(18736) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18736))))  severity failure;
	assert RAM(18737) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18737))))  severity failure;
	assert RAM(18738) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18738))))  severity failure;
	assert RAM(18739) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18739))))  severity failure;
	assert RAM(18740) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18740))))  severity failure;
	assert RAM(18741) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18741))))  severity failure;
	assert RAM(18742) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18742))))  severity failure;
	assert RAM(18743) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18743))))  severity failure;
	assert RAM(18744) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18744))))  severity failure;
	assert RAM(18745) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18745))))  severity failure;
	assert RAM(18746) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18746))))  severity failure;
	assert RAM(18747) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18747))))  severity failure;
	assert RAM(18748) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18748))))  severity failure;
	assert RAM(18749) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18749))))  severity failure;
	assert RAM(18750) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18750))))  severity failure;
	assert RAM(18751) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18751))))  severity failure;
	assert RAM(18752) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(18752))))  severity failure;
	assert RAM(18753) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18753))))  severity failure;
	assert RAM(18754) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18754))))  severity failure;
	assert RAM(18755) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18755))))  severity failure;
	assert RAM(18756) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18756))))  severity failure;
	assert RAM(18757) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(18757))))  severity failure;
	assert RAM(18758) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18758))))  severity failure;
	assert RAM(18759) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18759))))  severity failure;
	assert RAM(18760) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18760))))  severity failure;
	assert RAM(18761) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18761))))  severity failure;
	assert RAM(18762) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(18762))))  severity failure;
	assert RAM(18763) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18763))))  severity failure;
	assert RAM(18764) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18764))))  severity failure;
	assert RAM(18765) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18765))))  severity failure;
	assert RAM(18766) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18766))))  severity failure;
	assert RAM(18767) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18767))))  severity failure;
	assert RAM(18768) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18768))))  severity failure;
	assert RAM(18769) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18769))))  severity failure;
	assert RAM(18770) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18770))))  severity failure;
	assert RAM(18771) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(18771))))  severity failure;
	assert RAM(18772) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18772))))  severity failure;
	assert RAM(18773) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18773))))  severity failure;
	assert RAM(18774) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18774))))  severity failure;
	assert RAM(18775) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18775))))  severity failure;
	assert RAM(18776) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18776))))  severity failure;
	assert RAM(18777) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18777))))  severity failure;
	assert RAM(18778) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(18778))))  severity failure;
	assert RAM(18779) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18779))))  severity failure;
	assert RAM(18780) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18780))))  severity failure;
	assert RAM(18781) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(18781))))  severity failure;
	assert RAM(18782) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18782))))  severity failure;
	assert RAM(18783) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(18783))))  severity failure;
	assert RAM(18784) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18784))))  severity failure;
	assert RAM(18785) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18785))))  severity failure;
	assert RAM(18786) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18786))))  severity failure;
	assert RAM(18787) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18787))))  severity failure;
	assert RAM(18788) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18788))))  severity failure;
	assert RAM(18789) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18789))))  severity failure;
	assert RAM(18790) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18790))))  severity failure;
	assert RAM(18791) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18791))))  severity failure;
	assert RAM(18792) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18792))))  severity failure;
	assert RAM(18793) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18793))))  severity failure;
	assert RAM(18794) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18794))))  severity failure;
	assert RAM(18795) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(18795))))  severity failure;
	assert RAM(18796) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18796))))  severity failure;
	assert RAM(18797) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(18797))))  severity failure;
	assert RAM(18798) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18798))))  severity failure;
	assert RAM(18799) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(18799))))  severity failure;
	assert RAM(18800) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18800))))  severity failure;
	assert RAM(18801) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(18801))))  severity failure;
	assert RAM(18802) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18802))))  severity failure;
	assert RAM(18803) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18803))))  severity failure;
	assert RAM(18804) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18804))))  severity failure;
	assert RAM(18805) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(18805))))  severity failure;
	assert RAM(18806) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18806))))  severity failure;
	assert RAM(18807) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18807))))  severity failure;
	assert RAM(18808) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18808))))  severity failure;
	assert RAM(18809) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18809))))  severity failure;
	assert RAM(18810) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18810))))  severity failure;
	assert RAM(18811) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18811))))  severity failure;
	assert RAM(18812) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18812))))  severity failure;
	assert RAM(18813) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18813))))  severity failure;
	assert RAM(18814) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18814))))  severity failure;
	assert RAM(18815) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18815))))  severity failure;
	assert RAM(18816) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18816))))  severity failure;
	assert RAM(18817) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18817))))  severity failure;
	assert RAM(18818) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18818))))  severity failure;
	assert RAM(18819) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18819))))  severity failure;
	assert RAM(18820) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18820))))  severity failure;
	assert RAM(18821) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18821))))  severity failure;
	assert RAM(18822) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18822))))  severity failure;
	assert RAM(18823) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18823))))  severity failure;
	assert RAM(18824) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18824))))  severity failure;
	assert RAM(18825) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18825))))  severity failure;
	assert RAM(18826) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18826))))  severity failure;
	assert RAM(18827) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18827))))  severity failure;
	assert RAM(18828) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18828))))  severity failure;
	assert RAM(18829) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18829))))  severity failure;
	assert RAM(18830) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18830))))  severity failure;
	assert RAM(18831) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18831))))  severity failure;
	assert RAM(18832) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18832))))  severity failure;
	assert RAM(18833) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18833))))  severity failure;
	assert RAM(18834) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(18834))))  severity failure;
	assert RAM(18835) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18835))))  severity failure;
	assert RAM(18836) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18836))))  severity failure;
	assert RAM(18837) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18837))))  severity failure;
	assert RAM(18838) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18838))))  severity failure;
	assert RAM(18839) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18839))))  severity failure;
	assert RAM(18840) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18840))))  severity failure;
	assert RAM(18841) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18841))))  severity failure;
	assert RAM(18842) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(18842))))  severity failure;
	assert RAM(18843) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18843))))  severity failure;
	assert RAM(18844) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18844))))  severity failure;
	assert RAM(18845) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(18845))))  severity failure;
	assert RAM(18846) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18846))))  severity failure;
	assert RAM(18847) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18847))))  severity failure;
	assert RAM(18848) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18848))))  severity failure;
	assert RAM(18849) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18849))))  severity failure;
	assert RAM(18850) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(18850))))  severity failure;
	assert RAM(18851) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18851))))  severity failure;
	assert RAM(18852) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18852))))  severity failure;
	assert RAM(18853) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18853))))  severity failure;
	assert RAM(18854) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18854))))  severity failure;
	assert RAM(18855) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18855))))  severity failure;
	assert RAM(18856) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18856))))  severity failure;
	assert RAM(18857) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18857))))  severity failure;
	assert RAM(18858) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18858))))  severity failure;
	assert RAM(18859) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18859))))  severity failure;
	assert RAM(18860) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(18860))))  severity failure;
	assert RAM(18861) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(18861))))  severity failure;
	assert RAM(18862) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18862))))  severity failure;
	assert RAM(18863) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18863))))  severity failure;
	assert RAM(18864) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18864))))  severity failure;
	assert RAM(18865) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18865))))  severity failure;
	assert RAM(18866) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18866))))  severity failure;
	assert RAM(18867) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18867))))  severity failure;
	assert RAM(18868) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18868))))  severity failure;
	assert RAM(18869) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18869))))  severity failure;
	assert RAM(18870) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18870))))  severity failure;
	assert RAM(18871) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18871))))  severity failure;
	assert RAM(18872) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18872))))  severity failure;
	assert RAM(18873) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18873))))  severity failure;
	assert RAM(18874) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18874))))  severity failure;
	assert RAM(18875) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18875))))  severity failure;
	assert RAM(18876) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18876))))  severity failure;
	assert RAM(18877) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18877))))  severity failure;
	assert RAM(18878) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18878))))  severity failure;
	assert RAM(18879) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18879))))  severity failure;
	assert RAM(18880) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18880))))  severity failure;
	assert RAM(18881) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18881))))  severity failure;
	assert RAM(18882) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18882))))  severity failure;
	assert RAM(18883) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(18883))))  severity failure;
	assert RAM(18884) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18884))))  severity failure;
	assert RAM(18885) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18885))))  severity failure;
	assert RAM(18886) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18886))))  severity failure;
	assert RAM(18887) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18887))))  severity failure;
	assert RAM(18888) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18888))))  severity failure;
	assert RAM(18889) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18889))))  severity failure;
	assert RAM(18890) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18890))))  severity failure;
	assert RAM(18891) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18891))))  severity failure;
	assert RAM(18892) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18892))))  severity failure;
	assert RAM(18893) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18893))))  severity failure;
	assert RAM(18894) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18894))))  severity failure;
	assert RAM(18895) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18895))))  severity failure;
	assert RAM(18896) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18896))))  severity failure;
	assert RAM(18897) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18897))))  severity failure;
	assert RAM(18898) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18898))))  severity failure;
	assert RAM(18899) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18899))))  severity failure;
	assert RAM(18900) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18900))))  severity failure;
	assert RAM(18901) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18901))))  severity failure;
	assert RAM(18902) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(18902))))  severity failure;
	assert RAM(18903) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18903))))  severity failure;
	assert RAM(18904) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18904))))  severity failure;
	assert RAM(18905) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18905))))  severity failure;
	assert RAM(18906) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18906))))  severity failure;
	assert RAM(18907) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18907))))  severity failure;
	assert RAM(18908) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18908))))  severity failure;
	assert RAM(18909) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18909))))  severity failure;
	assert RAM(18910) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18910))))  severity failure;
	assert RAM(18911) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18911))))  severity failure;
	assert RAM(18912) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(18912))))  severity failure;
	assert RAM(18913) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18913))))  severity failure;
	assert RAM(18914) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18914))))  severity failure;
	assert RAM(18915) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18915))))  severity failure;
	assert RAM(18916) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18916))))  severity failure;
	assert RAM(18917) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18917))))  severity failure;
	assert RAM(18918) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(18918))))  severity failure;
	assert RAM(18919) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18919))))  severity failure;
	assert RAM(18920) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18920))))  severity failure;
	assert RAM(18921) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18921))))  severity failure;
	assert RAM(18922) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18922))))  severity failure;
	assert RAM(18923) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(18923))))  severity failure;
	assert RAM(18924) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18924))))  severity failure;
	assert RAM(18925) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18925))))  severity failure;
	assert RAM(18926) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18926))))  severity failure;
	assert RAM(18927) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18927))))  severity failure;
	assert RAM(18928) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18928))))  severity failure;
	assert RAM(18929) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18929))))  severity failure;
	assert RAM(18930) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18930))))  severity failure;
	assert RAM(18931) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18931))))  severity failure;
	assert RAM(18932) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18932))))  severity failure;
	assert RAM(18933) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(18933))))  severity failure;
	assert RAM(18934) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18934))))  severity failure;
	assert RAM(18935) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18935))))  severity failure;
	assert RAM(18936) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18936))))  severity failure;
	assert RAM(18937) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18937))))  severity failure;
	assert RAM(18938) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18938))))  severity failure;
	assert RAM(18939) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18939))))  severity failure;
	assert RAM(18940) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18940))))  severity failure;
	assert RAM(18941) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(18941))))  severity failure;
	assert RAM(18942) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(18942))))  severity failure;
	assert RAM(18943) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18943))))  severity failure;
	assert RAM(18944) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18944))))  severity failure;
	assert RAM(18945) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18945))))  severity failure;
	assert RAM(18946) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18946))))  severity failure;
	assert RAM(18947) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(18947))))  severity failure;
	assert RAM(18948) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18948))))  severity failure;
	assert RAM(18949) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18949))))  severity failure;
	assert RAM(18950) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18950))))  severity failure;
	assert RAM(18951) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18951))))  severity failure;
	assert RAM(18952) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18952))))  severity failure;
	assert RAM(18953) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18953))))  severity failure;
	assert RAM(18954) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18954))))  severity failure;
	assert RAM(18955) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18955))))  severity failure;
	assert RAM(18956) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18956))))  severity failure;
	assert RAM(18957) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18957))))  severity failure;
	assert RAM(18958) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18958))))  severity failure;
	assert RAM(18959) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18959))))  severity failure;
	assert RAM(18960) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(18960))))  severity failure;
	assert RAM(18961) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18961))))  severity failure;
	assert RAM(18962) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18962))))  severity failure;
	assert RAM(18963) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(18963))))  severity failure;
	assert RAM(18964) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18964))))  severity failure;
	assert RAM(18965) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18965))))  severity failure;
	assert RAM(18966) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18966))))  severity failure;
	assert RAM(18967) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18967))))  severity failure;
	assert RAM(18968) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18968))))  severity failure;
	assert RAM(18969) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18969))))  severity failure;
	assert RAM(18970) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18970))))  severity failure;
	assert RAM(18971) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18971))))  severity failure;
	assert RAM(18972) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18972))))  severity failure;
	assert RAM(18973) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18973))))  severity failure;
	assert RAM(18974) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18974))))  severity failure;
	assert RAM(18975) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18975))))  severity failure;
	assert RAM(18976) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18976))))  severity failure;
	assert RAM(18977) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18977))))  severity failure;
	assert RAM(18978) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18978))))  severity failure;
	assert RAM(18979) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18979))))  severity failure;
	assert RAM(18980) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18980))))  severity failure;
	assert RAM(18981) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18981))))  severity failure;
	assert RAM(18982) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(18982))))  severity failure;
	assert RAM(18983) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18983))))  severity failure;
	assert RAM(18984) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18984))))  severity failure;
	assert RAM(18985) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18985))))  severity failure;
	assert RAM(18986) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18986))))  severity failure;
	assert RAM(18987) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18987))))  severity failure;
	assert RAM(18988) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18988))))  severity failure;
	assert RAM(18989) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18989))))  severity failure;
	assert RAM(18990) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18990))))  severity failure;
	assert RAM(18991) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18991))))  severity failure;
	assert RAM(18992) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18992))))  severity failure;
	assert RAM(18993) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18993))))  severity failure;
	assert RAM(18994) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18994))))  severity failure;
	assert RAM(18995) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18995))))  severity failure;
	assert RAM(18996) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18996))))  severity failure;
	assert RAM(18997) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18997))))  severity failure;
	assert RAM(18998) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18998))))  severity failure;
	assert RAM(18999) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18999))))  severity failure;
	assert RAM(19000) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(19000))))  severity failure;
	assert RAM(19001) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19001))))  severity failure;
	assert RAM(19002) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(19002))))  severity failure;
	assert RAM(19003) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19003))))  severity failure;
	assert RAM(19004) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19004))))  severity failure;
	assert RAM(19005) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19005))))  severity failure;
	assert RAM(19006) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19006))))  severity failure;
	assert RAM(19007) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19007))))  severity failure;
	assert RAM(19008) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19008))))  severity failure;
	assert RAM(19009) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19009))))  severity failure;
	assert RAM(19010) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19010))))  severity failure;
	assert RAM(19011) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19011))))  severity failure;
	assert RAM(19012) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19012))))  severity failure;
	assert RAM(19013) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(19013))))  severity failure;
	assert RAM(19014) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19014))))  severity failure;
	assert RAM(19015) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19015))))  severity failure;
	assert RAM(19016) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19016))))  severity failure;
	assert RAM(19017) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19017))))  severity failure;
	assert RAM(19018) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19018))))  severity failure;
	assert RAM(19019) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19019))))  severity failure;
	assert RAM(19020) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19020))))  severity failure;
	assert RAM(19021) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19021))))  severity failure;
	assert RAM(19022) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(19022))))  severity failure;
	assert RAM(19023) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19023))))  severity failure;
	assert RAM(19024) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19024))))  severity failure;
	assert RAM(19025) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19025))))  severity failure;
	assert RAM(19026) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19026))))  severity failure;
	assert RAM(19027) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19027))))  severity failure;
	assert RAM(19028) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19028))))  severity failure;
	assert RAM(19029) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19029))))  severity failure;
	assert RAM(19030) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19030))))  severity failure;
	assert RAM(19031) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19031))))  severity failure;
	assert RAM(19032) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19032))))  severity failure;
	assert RAM(19033) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19033))))  severity failure;
	assert RAM(19034) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19034))))  severity failure;
	assert RAM(19035) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19035))))  severity failure;
	assert RAM(19036) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(19036))))  severity failure;
	assert RAM(19037) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19037))))  severity failure;
	assert RAM(19038) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19038))))  severity failure;
	assert RAM(19039) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19039))))  severity failure;
	assert RAM(19040) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19040))))  severity failure;
	assert RAM(19041) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19041))))  severity failure;
	assert RAM(19042) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19042))))  severity failure;
	assert RAM(19043) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19043))))  severity failure;
	assert RAM(19044) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19044))))  severity failure;
	assert RAM(19045) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19045))))  severity failure;
	assert RAM(19046) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(19046))))  severity failure;
	assert RAM(19047) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19047))))  severity failure;
	assert RAM(19048) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19048))))  severity failure;
	assert RAM(19049) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19049))))  severity failure;
	assert RAM(19050) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19050))))  severity failure;
	assert RAM(19051) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(19051))))  severity failure;
	assert RAM(19052) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19052))))  severity failure;
	assert RAM(19053) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19053))))  severity failure;
	assert RAM(19054) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19054))))  severity failure;
	assert RAM(19055) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19055))))  severity failure;
	assert RAM(19056) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19056))))  severity failure;
	assert RAM(19057) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19057))))  severity failure;
	assert RAM(19058) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19058))))  severity failure;
	assert RAM(19059) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19059))))  severity failure;
	assert RAM(19060) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19060))))  severity failure;
	assert RAM(19061) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19061))))  severity failure;
	assert RAM(19062) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19062))))  severity failure;
	assert RAM(19063) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19063))))  severity failure;
	assert RAM(19064) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(19064))))  severity failure;
	assert RAM(19065) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19065))))  severity failure;
	assert RAM(19066) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19066))))  severity failure;
	assert RAM(19067) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(19067))))  severity failure;
	assert RAM(19068) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19068))))  severity failure;
	assert RAM(19069) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19069))))  severity failure;
	assert RAM(19070) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19070))))  severity failure;
	assert RAM(19071) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19071))))  severity failure;
	assert RAM(19072) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(19072))))  severity failure;
	assert RAM(19073) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19073))))  severity failure;
	assert RAM(19074) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19074))))  severity failure;
	assert RAM(19075) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(19075))))  severity failure;
	assert RAM(19076) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19076))))  severity failure;
	assert RAM(19077) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19077))))  severity failure;
	assert RAM(19078) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19078))))  severity failure;
	assert RAM(19079) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19079))))  severity failure;
	assert RAM(19080) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19080))))  severity failure;
	assert RAM(19081) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19081))))  severity failure;
	assert RAM(19082) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19082))))  severity failure;
	assert RAM(19083) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19083))))  severity failure;
	assert RAM(19084) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19084))))  severity failure;
	assert RAM(19085) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19085))))  severity failure;
	assert RAM(19086) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19086))))  severity failure;
	assert RAM(19087) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19087))))  severity failure;
	assert RAM(19088) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19088))))  severity failure;
	assert RAM(19089) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19089))))  severity failure;
	assert RAM(19090) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19090))))  severity failure;
	assert RAM(19091) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19091))))  severity failure;
	assert RAM(19092) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(19092))))  severity failure;
	assert RAM(19093) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19093))))  severity failure;
	assert RAM(19094) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19094))))  severity failure;
	assert RAM(19095) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19095))))  severity failure;
	assert RAM(19096) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19096))))  severity failure;
	assert RAM(19097) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(19097))))  severity failure;
	assert RAM(19098) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(19098))))  severity failure;
	assert RAM(19099) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19099))))  severity failure;
	assert RAM(19100) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19100))))  severity failure;
	assert RAM(19101) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19101))))  severity failure;
	assert RAM(19102) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19102))))  severity failure;
	assert RAM(19103) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19103))))  severity failure;
	assert RAM(19104) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19104))))  severity failure;
	assert RAM(19105) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19105))))  severity failure;
	assert RAM(19106) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19106))))  severity failure;
	assert RAM(19107) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19107))))  severity failure;
	assert RAM(19108) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19108))))  severity failure;
	assert RAM(19109) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19109))))  severity failure;
	assert RAM(19110) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19110))))  severity failure;
	assert RAM(19111) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(19111))))  severity failure;
	assert RAM(19112) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19112))))  severity failure;
	assert RAM(19113) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(19113))))  severity failure;
	assert RAM(19114) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19114))))  severity failure;
	assert RAM(19115) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19115))))  severity failure;
	assert RAM(19116) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19116))))  severity failure;
	assert RAM(19117) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(19117))))  severity failure;
	assert RAM(19118) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19118))))  severity failure;
	assert RAM(19119) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(19119))))  severity failure;
	assert RAM(19120) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19120))))  severity failure;
	assert RAM(19121) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19121))))  severity failure;
	assert RAM(19122) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19122))))  severity failure;
	assert RAM(19123) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19123))))  severity failure;
	assert RAM(19124) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19124))))  severity failure;
	assert RAM(19125) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(19125))))  severity failure;
	assert RAM(19126) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19126))))  severity failure;
	assert RAM(19127) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19127))))  severity failure;
	assert RAM(19128) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19128))))  severity failure;
	assert RAM(19129) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19129))))  severity failure;
	assert RAM(19130) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19130))))  severity failure;
	assert RAM(19131) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19131))))  severity failure;
	assert RAM(19132) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19132))))  severity failure;
	assert RAM(19133) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19133))))  severity failure;
	assert RAM(19134) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19134))))  severity failure;
	assert RAM(19135) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(19135))))  severity failure;
	assert RAM(19136) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(19136))))  severity failure;
	assert RAM(19137) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19137))))  severity failure;
	assert RAM(19138) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19138))))  severity failure;
	assert RAM(19139) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19139))))  severity failure;
	assert RAM(19140) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19140))))  severity failure;
	assert RAM(19141) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19141))))  severity failure;
	assert RAM(19142) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19142))))  severity failure;
	assert RAM(19143) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19143))))  severity failure;
	assert RAM(19144) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19144))))  severity failure;
	assert RAM(19145) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19145))))  severity failure;
	assert RAM(19146) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19146))))  severity failure;
	assert RAM(19147) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19147))))  severity failure;
	assert RAM(19148) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19148))))  severity failure;
	assert RAM(19149) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19149))))  severity failure;
	assert RAM(19150) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19150))))  severity failure;
	assert RAM(19151) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19151))))  severity failure;
	assert RAM(19152) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19152))))  severity failure;
	assert RAM(19153) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19153))))  severity failure;
	assert RAM(19154) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19154))))  severity failure;
	assert RAM(19155) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19155))))  severity failure;
	assert RAM(19156) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19156))))  severity failure;
	assert RAM(19157) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19157))))  severity failure;
	assert RAM(19158) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19158))))  severity failure;
	assert RAM(19159) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19159))))  severity failure;
	assert RAM(19160) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19160))))  severity failure;
	assert RAM(19161) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19161))))  severity failure;
	assert RAM(19162) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19162))))  severity failure;
	assert RAM(19163) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19163))))  severity failure;
	assert RAM(19164) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(19164))))  severity failure;
	assert RAM(19165) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19165))))  severity failure;
	assert RAM(19166) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19166))))  severity failure;
	assert RAM(19167) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19167))))  severity failure;
	assert RAM(19168) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19168))))  severity failure;
	assert RAM(19169) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19169))))  severity failure;
	assert RAM(19170) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19170))))  severity failure;
	assert RAM(19171) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19171))))  severity failure;
	assert RAM(19172) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19172))))  severity failure;
	assert RAM(19173) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19173))))  severity failure;
	assert RAM(19174) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19174))))  severity failure;
	assert RAM(19175) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19175))))  severity failure;
	assert RAM(19176) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19176))))  severity failure;
	assert RAM(19177) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19177))))  severity failure;
	assert RAM(19178) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19178))))  severity failure;
	assert RAM(19179) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19179))))  severity failure;
	assert RAM(19180) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19180))))  severity failure;
	assert RAM(19181) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19181))))  severity failure;
	assert RAM(19182) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19182))))  severity failure;
	assert RAM(19183) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(19183))))  severity failure;
	assert RAM(19184) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19184))))  severity failure;
	assert RAM(19185) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19185))))  severity failure;
	assert RAM(19186) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19186))))  severity failure;
	assert RAM(19187) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19187))))  severity failure;
	assert RAM(19188) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(19188))))  severity failure;
	assert RAM(19189) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(19189))))  severity failure;
	assert RAM(19190) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19190))))  severity failure;
	assert RAM(19191) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19191))))  severity failure;
	assert RAM(19192) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19192))))  severity failure;
	assert RAM(19193) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19193))))  severity failure;
	assert RAM(19194) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19194))))  severity failure;
	assert RAM(19195) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19195))))  severity failure;
	assert RAM(19196) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19196))))  severity failure;
	assert RAM(19197) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19197))))  severity failure;
	assert RAM(19198) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(19198))))  severity failure;
	assert RAM(19199) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19199))))  severity failure;
	assert RAM(19200) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19200))))  severity failure;
	assert RAM(19201) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19201))))  severity failure;
	assert RAM(19202) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19202))))  severity failure;
	assert RAM(19203) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19203))))  severity failure;
	assert RAM(19204) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19204))))  severity failure;
	assert RAM(19205) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19205))))  severity failure;
	assert RAM(19206) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19206))))  severity failure;
	assert RAM(19207) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(19207))))  severity failure;
	assert RAM(19208) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19208))))  severity failure;
	assert RAM(19209) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(19209))))  severity failure;
	assert RAM(19210) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(19210))))  severity failure;
	assert RAM(19211) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19211))))  severity failure;
	assert RAM(19212) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(19212))))  severity failure;
	assert RAM(19213) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19213))))  severity failure;
	assert RAM(19214) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19214))))  severity failure;
	assert RAM(19215) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19215))))  severity failure;
	assert RAM(19216) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19216))))  severity failure;
	assert RAM(19217) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(19217))))  severity failure;
	assert RAM(19218) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19218))))  severity failure;
	assert RAM(19219) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19219))))  severity failure;
	assert RAM(19220) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19220))))  severity failure;
	assert RAM(19221) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19221))))  severity failure;
	assert RAM(19222) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19222))))  severity failure;
	assert RAM(19223) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19223))))  severity failure;
	assert RAM(19224) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19224))))  severity failure;
	assert RAM(19225) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19225))))  severity failure;
	assert RAM(19226) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19226))))  severity failure;
	assert RAM(19227) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19227))))  severity failure;
	assert RAM(19228) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19228))))  severity failure;
	assert RAM(19229) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19229))))  severity failure;
	assert RAM(19230) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19230))))  severity failure;
	assert RAM(19231) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19231))))  severity failure;
	assert RAM(19232) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19232))))  severity failure;
	assert RAM(19233) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19233))))  severity failure;
	assert RAM(19234) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(19234))))  severity failure;
	assert RAM(19235) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19235))))  severity failure;
	assert RAM(19236) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(19236))))  severity failure;
	assert RAM(19237) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19237))))  severity failure;
	assert RAM(19238) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19238))))  severity failure;
	assert RAM(19239) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19239))))  severity failure;
	assert RAM(19240) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19240))))  severity failure;
	assert RAM(19241) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19241))))  severity failure;
	assert RAM(19242) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19242))))  severity failure;
	assert RAM(19243) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(19243))))  severity failure;
	assert RAM(19244) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19244))))  severity failure;
	assert RAM(19245) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19245))))  severity failure;
	assert RAM(19246) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19246))))  severity failure;
	assert RAM(19247) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19247))))  severity failure;
	assert RAM(19248) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19248))))  severity failure;
	assert RAM(19249) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(19249))))  severity failure;
	assert RAM(19250) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19250))))  severity failure;
	assert RAM(19251) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19251))))  severity failure;
	assert RAM(19252) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19252))))  severity failure;
	assert RAM(19253) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19253))))  severity failure;
	assert RAM(19254) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19254))))  severity failure;
	assert RAM(19255) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19255))))  severity failure;
	assert RAM(19256) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19256))))  severity failure;
	assert RAM(19257) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19257))))  severity failure;
	assert RAM(19258) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19258))))  severity failure;
	assert RAM(19259) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19259))))  severity failure;
	assert RAM(19260) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19260))))  severity failure;
	assert RAM(19261) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19261))))  severity failure;
	assert RAM(19262) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19262))))  severity failure;
	assert RAM(19263) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19263))))  severity failure;
	assert RAM(19264) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19264))))  severity failure;
	assert RAM(19265) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19265))))  severity failure;
	assert RAM(19266) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(19266))))  severity failure;
	assert RAM(19267) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19267))))  severity failure;
	assert RAM(19268) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19268))))  severity failure;
	assert RAM(19269) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(19269))))  severity failure;
	assert RAM(19270) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19270))))  severity failure;
	assert RAM(19271) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19271))))  severity failure;
	assert RAM(19272) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19272))))  severity failure;
	assert RAM(19273) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(19273))))  severity failure;
	assert RAM(19274) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19274))))  severity failure;
	assert RAM(19275) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19275))))  severity failure;
	assert RAM(19276) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19276))))  severity failure;
	assert RAM(19277) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19277))))  severity failure;
	assert RAM(19278) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19278))))  severity failure;
	assert RAM(19279) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19279))))  severity failure;
	assert RAM(19280) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19280))))  severity failure;
	assert RAM(19281) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19281))))  severity failure;
	assert RAM(19282) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19282))))  severity failure;
	assert RAM(19283) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19283))))  severity failure;
	assert RAM(19284) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19284))))  severity failure;
	assert RAM(19285) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(19285))))  severity failure;
	assert RAM(19286) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19286))))  severity failure;
	assert RAM(19287) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19287))))  severity failure;
	assert RAM(19288) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19288))))  severity failure;
	assert RAM(19289) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(19289))))  severity failure;
	assert RAM(19290) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19290))))  severity failure;
	assert RAM(19291) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19291))))  severity failure;
	assert RAM(19292) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19292))))  severity failure;
	assert RAM(19293) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(19293))))  severity failure;
	assert RAM(19294) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19294))))  severity failure;
	assert RAM(19295) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(19295))))  severity failure;
	assert RAM(19296) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19296))))  severity failure;
	assert RAM(19297) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19297))))  severity failure;
	assert RAM(19298) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19298))))  severity failure;
	assert RAM(19299) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19299))))  severity failure;
	assert RAM(19300) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19300))))  severity failure;
	assert RAM(19301) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19301))))  severity failure;
	assert RAM(19302) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19302))))  severity failure;
	assert RAM(19303) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19303))))  severity failure;
	assert RAM(19304) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19304))))  severity failure;
	assert RAM(19305) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19305))))  severity failure;
	assert RAM(19306) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(19306))))  severity failure;
	assert RAM(19307) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19307))))  severity failure;
	assert RAM(19308) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19308))))  severity failure;
	assert RAM(19309) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19309))))  severity failure;
	assert RAM(19310) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(19310))))  severity failure;
	assert RAM(19311) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(19311))))  severity failure;
	assert RAM(19312) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19312))))  severity failure;
	assert RAM(19313) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19313))))  severity failure;
	assert RAM(19314) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19314))))  severity failure;
	assert RAM(19315) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19315))))  severity failure;
	assert RAM(19316) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19316))))  severity failure;
	assert RAM(19317) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19317))))  severity failure;
	assert RAM(19318) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19318))))  severity failure;
	assert RAM(19319) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19319))))  severity failure;
	assert RAM(19320) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19320))))  severity failure;
	assert RAM(19321) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(19321))))  severity failure;
	assert RAM(19322) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19322))))  severity failure;
	assert RAM(19323) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19323))))  severity failure;
	assert RAM(19324) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19324))))  severity failure;
	assert RAM(19325) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19325))))  severity failure;
	assert RAM(19326) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19326))))  severity failure;
	assert RAM(19327) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19327))))  severity failure;
	assert RAM(19328) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19328))))  severity failure;
	assert RAM(19329) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19329))))  severity failure;
	assert RAM(19330) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19330))))  severity failure;
	assert RAM(19331) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19331))))  severity failure;
	assert RAM(19332) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19332))))  severity failure;
	assert RAM(19333) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(19333))))  severity failure;
	assert RAM(19334) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19334))))  severity failure;
	assert RAM(19335) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19335))))  severity failure;
	assert RAM(19336) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19336))))  severity failure;
	assert RAM(19337) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19337))))  severity failure;
	assert RAM(19338) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19338))))  severity failure;
	assert RAM(19339) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19339))))  severity failure;
	assert RAM(19340) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(19340))))  severity failure;
	assert RAM(19341) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19341))))  severity failure;
	assert RAM(19342) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19342))))  severity failure;
	assert RAM(19343) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19343))))  severity failure;
	assert RAM(19344) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19344))))  severity failure;
	assert RAM(19345) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19345))))  severity failure;
	assert RAM(19346) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19346))))  severity failure;
	assert RAM(19347) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19347))))  severity failure;
	assert RAM(19348) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19348))))  severity failure;
	assert RAM(19349) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19349))))  severity failure;
	assert RAM(19350) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19350))))  severity failure;
	assert RAM(19351) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19351))))  severity failure;
	assert RAM(19352) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(19352))))  severity failure;
	assert RAM(19353) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(19353))))  severity failure;
	assert RAM(19354) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(19354))))  severity failure;
	assert RAM(19355) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19355))))  severity failure;
	assert RAM(19356) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19356))))  severity failure;
	assert RAM(19357) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(19357))))  severity failure;
	assert RAM(19358) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19358))))  severity failure;
	assert RAM(19359) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19359))))  severity failure;
	assert RAM(19360) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19360))))  severity failure;
	assert RAM(19361) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19361))))  severity failure;
	assert RAM(19362) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19362))))  severity failure;
	assert RAM(19363) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19363))))  severity failure;
	assert RAM(19364) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19364))))  severity failure;
	assert RAM(19365) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(19365))))  severity failure;
	assert RAM(19366) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19366))))  severity failure;
	assert RAM(19367) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19367))))  severity failure;
	assert RAM(19368) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19368))))  severity failure;
	assert RAM(19369) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19369))))  severity failure;
	assert RAM(19370) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19370))))  severity failure;
	assert RAM(19371) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19371))))  severity failure;
	assert RAM(19372) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19372))))  severity failure;
	assert RAM(19373) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(19373))))  severity failure;
	assert RAM(19374) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19374))))  severity failure;
	assert RAM(19375) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19375))))  severity failure;
	assert RAM(19376) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19376))))  severity failure;
	assert RAM(19377) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(19377))))  severity failure;
	assert RAM(19378) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19378))))  severity failure;
	assert RAM(19379) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(19379))))  severity failure;
	assert RAM(19380) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19380))))  severity failure;
	assert RAM(19381) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(19381))))  severity failure;
	assert RAM(19382) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19382))))  severity failure;
	assert RAM(19383) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19383))))  severity failure;
	assert RAM(19384) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19384))))  severity failure;
	assert RAM(19385) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19385))))  severity failure;
	assert RAM(19386) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19386))))  severity failure;
	assert RAM(19387) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19387))))  severity failure;
	assert RAM(19388) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19388))))  severity failure;
	assert RAM(19389) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19389))))  severity failure;
	assert RAM(19390) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19390))))  severity failure;
	assert RAM(19391) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(19391))))  severity failure;
	assert RAM(19392) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19392))))  severity failure;
	assert RAM(19393) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19393))))  severity failure;
	assert RAM(19394) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19394))))  severity failure;
	assert RAM(19395) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19395))))  severity failure;
	assert RAM(19396) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19396))))  severity failure;
	assert RAM(19397) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19397))))  severity failure;
	assert RAM(19398) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19398))))  severity failure;
	assert RAM(19399) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19399))))  severity failure;
	assert RAM(19400) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19400))))  severity failure;
	assert RAM(19401) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19401))))  severity failure;
	assert RAM(19402) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19402))))  severity failure;
	assert RAM(19403) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19403))))  severity failure;
	assert RAM(19404) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19404))))  severity failure;
	assert RAM(19405) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19405))))  severity failure;
	assert RAM(19406) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19406))))  severity failure;
	assert RAM(19407) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19407))))  severity failure;
	assert RAM(19408) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(19408))))  severity failure;
	assert RAM(19409) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19409))))  severity failure;
	assert RAM(19410) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19410))))  severity failure;
	assert RAM(19411) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19411))))  severity failure;
	assert RAM(19412) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19412))))  severity failure;
	assert RAM(19413) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19413))))  severity failure;
	assert RAM(19414) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19414))))  severity failure;
	assert RAM(19415) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19415))))  severity failure;
	assert RAM(19416) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19416))))  severity failure;
	assert RAM(19417) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19417))))  severity failure;
	assert RAM(19418) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19418))))  severity failure;
	assert RAM(19419) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19419))))  severity failure;
	assert RAM(19420) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19420))))  severity failure;
	assert RAM(19421) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19421))))  severity failure;
	assert RAM(19422) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19422))))  severity failure;
	assert RAM(19423) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19423))))  severity failure;
	assert RAM(19424) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19424))))  severity failure;
	assert RAM(19425) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19425))))  severity failure;
	assert RAM(19426) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19426))))  severity failure;
	assert RAM(19427) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19427))))  severity failure;
	assert RAM(19428) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19428))))  severity failure;
	assert RAM(19429) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19429))))  severity failure;
	assert RAM(19430) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19430))))  severity failure;
	assert RAM(19431) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19431))))  severity failure;
	assert RAM(19432) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19432))))  severity failure;
	assert RAM(19433) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19433))))  severity failure;
	assert RAM(19434) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(19434))))  severity failure;
	assert RAM(19435) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(19435))))  severity failure;
	assert RAM(19436) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19436))))  severity failure;
	assert RAM(19437) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19437))))  severity failure;
	assert RAM(19438) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(19438))))  severity failure;
	assert RAM(19439) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19439))))  severity failure;
	assert RAM(19440) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19440))))  severity failure;
	assert RAM(19441) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19441))))  severity failure;
	assert RAM(19442) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19442))))  severity failure;
	assert RAM(19443) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19443))))  severity failure;
	assert RAM(19444) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19444))))  severity failure;
	assert RAM(19445) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19445))))  severity failure;
	assert RAM(19446) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19446))))  severity failure;
	assert RAM(19447) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19447))))  severity failure;
	assert RAM(19448) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19448))))  severity failure;
	assert RAM(19449) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19449))))  severity failure;
	assert RAM(19450) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19450))))  severity failure;
	assert RAM(19451) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19451))))  severity failure;
	assert RAM(19452) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19452))))  severity failure;
	assert RAM(19453) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19453))))  severity failure;
	assert RAM(19454) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19454))))  severity failure;
	assert RAM(19455) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19455))))  severity failure;
	assert RAM(19456) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19456))))  severity failure;
	assert RAM(19457) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19457))))  severity failure;
	assert RAM(19458) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19458))))  severity failure;
	assert RAM(19459) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19459))))  severity failure;
	assert RAM(19460) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19460))))  severity failure;
	assert RAM(19461) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19461))))  severity failure;
	assert RAM(19462) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19462))))  severity failure;
	assert RAM(19463) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(19463))))  severity failure;
	assert RAM(19464) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19464))))  severity failure;
	assert RAM(19465) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19465))))  severity failure;
	assert RAM(19466) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19466))))  severity failure;
	assert RAM(19467) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19467))))  severity failure;
	assert RAM(19468) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19468))))  severity failure;
	assert RAM(19469) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19469))))  severity failure;
	assert RAM(19470) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19470))))  severity failure;
	assert RAM(19471) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19471))))  severity failure;
	assert RAM(19472) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19472))))  severity failure;
	assert RAM(19473) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19473))))  severity failure;
	assert RAM(19474) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19474))))  severity failure;
	assert RAM(19475) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19475))))  severity failure;
	assert RAM(19476) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19476))))  severity failure;
	assert RAM(19477) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19477))))  severity failure;
	assert RAM(19478) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19478))))  severity failure;
	assert RAM(19479) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(19479))))  severity failure;
	assert RAM(19480) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19480))))  severity failure;
	assert RAM(19481) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19481))))  severity failure;
	assert RAM(19482) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19482))))  severity failure;
	assert RAM(19483) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19483))))  severity failure;
	assert RAM(19484) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19484))))  severity failure;
	assert RAM(19485) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19485))))  severity failure;
	assert RAM(19486) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19486))))  severity failure;
	assert RAM(19487) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19487))))  severity failure;
	assert RAM(19488) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19488))))  severity failure;
	assert RAM(19489) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(19489))))  severity failure;
	assert RAM(19490) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19490))))  severity failure;
	assert RAM(19491) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19491))))  severity failure;
	assert RAM(19492) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19492))))  severity failure;
	assert RAM(19493) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19493))))  severity failure;
	assert RAM(19494) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19494))))  severity failure;
	assert RAM(19495) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19495))))  severity failure;
	assert RAM(19496) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19496))))  severity failure;
	assert RAM(19497) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19497))))  severity failure;
	assert RAM(19498) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19498))))  severity failure;
	assert RAM(19499) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19499))))  severity failure;
	assert RAM(19500) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19500))))  severity failure;
	assert RAM(19501) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(19501))))  severity failure;
	assert RAM(19502) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(19502))))  severity failure;
	assert RAM(19503) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19503))))  severity failure;
	assert RAM(19504) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19504))))  severity failure;
	assert RAM(19505) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19505))))  severity failure;
	assert RAM(19506) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19506))))  severity failure;
	assert RAM(19507) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19507))))  severity failure;
	assert RAM(19508) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19508))))  severity failure;
	assert RAM(19509) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19509))))  severity failure;
	assert RAM(19510) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19510))))  severity failure;
	assert RAM(19511) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19511))))  severity failure;
	assert RAM(19512) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19512))))  severity failure;
	assert RAM(19513) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19513))))  severity failure;
	assert RAM(19514) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19514))))  severity failure;
	assert RAM(19515) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(19515))))  severity failure;
	assert RAM(19516) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19516))))  severity failure;
	assert RAM(19517) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19517))))  severity failure;
	assert RAM(19518) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19518))))  severity failure;
	assert RAM(19519) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19519))))  severity failure;
	assert RAM(19520) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19520))))  severity failure;
	assert RAM(19521) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19521))))  severity failure;
	assert RAM(19522) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19522))))  severity failure;
	assert RAM(19523) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19523))))  severity failure;
	assert RAM(19524) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19524))))  severity failure;
	assert RAM(19525) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19525))))  severity failure;
	assert RAM(19526) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19526))))  severity failure;
	assert RAM(19527) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19527))))  severity failure;
	assert RAM(19528) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19528))))  severity failure;
	assert RAM(19529) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19529))))  severity failure;
	assert RAM(19530) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19530))))  severity failure;
	assert RAM(19531) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19531))))  severity failure;
	assert RAM(19532) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(19532))))  severity failure;
	assert RAM(19533) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19533))))  severity failure;
	assert RAM(19534) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19534))))  severity failure;
	assert RAM(19535) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19535))))  severity failure;
	assert RAM(19536) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19536))))  severity failure;
	assert RAM(19537) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19537))))  severity failure;
	assert RAM(19538) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19538))))  severity failure;
	assert RAM(19539) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19539))))  severity failure;
	assert RAM(19540) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19540))))  severity failure;
	assert RAM(19541) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19541))))  severity failure;
	assert RAM(19542) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19542))))  severity failure;
	assert RAM(19543) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19543))))  severity failure;
	assert RAM(19544) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19544))))  severity failure;
	assert RAM(19545) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19545))))  severity failure;
	assert RAM(19546) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19546))))  severity failure;
	assert RAM(19547) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19547))))  severity failure;
	assert RAM(19548) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19548))))  severity failure;
	assert RAM(19549) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19549))))  severity failure;
	assert RAM(19550) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(19550))))  severity failure;
	assert RAM(19551) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19551))))  severity failure;
	assert RAM(19552) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19552))))  severity failure;
	assert RAM(19553) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19553))))  severity failure;
	assert RAM(19554) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19554))))  severity failure;
	assert RAM(19555) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19555))))  severity failure;
	assert RAM(19556) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19556))))  severity failure;
	assert RAM(19557) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19557))))  severity failure;
	assert RAM(19558) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19558))))  severity failure;
	assert RAM(19559) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(19559))))  severity failure;
	assert RAM(19560) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19560))))  severity failure;
	assert RAM(19561) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19561))))  severity failure;
	assert RAM(19562) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19562))))  severity failure;
	assert RAM(19563) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(19563))))  severity failure;
	assert RAM(19564) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19564))))  severity failure;
	assert RAM(19565) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19565))))  severity failure;
	assert RAM(19566) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19566))))  severity failure;
	assert RAM(19567) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19567))))  severity failure;
	assert RAM(19568) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19568))))  severity failure;
	assert RAM(19569) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(19569))))  severity failure;
	assert RAM(19570) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19570))))  severity failure;
	assert RAM(19571) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19571))))  severity failure;
	assert RAM(19572) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19572))))  severity failure;
	assert RAM(19573) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(19573))))  severity failure;
	assert RAM(19574) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19574))))  severity failure;
	assert RAM(19575) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19575))))  severity failure;
	assert RAM(19576) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19576))))  severity failure;
	assert RAM(19577) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19577))))  severity failure;
	assert RAM(19578) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19578))))  severity failure;
	assert RAM(19579) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19579))))  severity failure;
	assert RAM(19580) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19580))))  severity failure;
	assert RAM(19581) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19581))))  severity failure;
	assert RAM(19582) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19582))))  severity failure;
	assert RAM(19583) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19583))))  severity failure;
	assert RAM(19584) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19584))))  severity failure;
	assert RAM(19585) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19585))))  severity failure;
	assert RAM(19586) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19586))))  severity failure;
	assert RAM(19587) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19587))))  severity failure;
	assert RAM(19588) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19588))))  severity failure;
	assert RAM(19589) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19589))))  severity failure;
	assert RAM(19590) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19590))))  severity failure;
	assert RAM(19591) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19591))))  severity failure;
	assert RAM(19592) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19592))))  severity failure;
	assert RAM(19593) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19593))))  severity failure;
	assert RAM(19594) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19594))))  severity failure;
	assert RAM(19595) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19595))))  severity failure;
	assert RAM(19596) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19596))))  severity failure;
	assert RAM(19597) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19597))))  severity failure;
	assert RAM(19598) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19598))))  severity failure;
	assert RAM(19599) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19599))))  severity failure;
	assert RAM(19600) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19600))))  severity failure;
	assert RAM(19601) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19601))))  severity failure;
	assert RAM(19602) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19602))))  severity failure;
	assert RAM(19603) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19603))))  severity failure;
	assert RAM(19604) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19604))))  severity failure;
	assert RAM(19605) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19605))))  severity failure;
	assert RAM(19606) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19606))))  severity failure;
	assert RAM(19607) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19607))))  severity failure;
	assert RAM(19608) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19608))))  severity failure;
	assert RAM(19609) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19609))))  severity failure;
	assert RAM(19610) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19610))))  severity failure;
	assert RAM(19611) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19611))))  severity failure;
	assert RAM(19612) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19612))))  severity failure;
	assert RAM(19613) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19613))))  severity failure;
	assert RAM(19614) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19614))))  severity failure;
	assert RAM(19615) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19615))))  severity failure;
	assert RAM(19616) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19616))))  severity failure;
	assert RAM(19617) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19617))))  severity failure;
	assert RAM(19618) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19618))))  severity failure;
	assert RAM(19619) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19619))))  severity failure;
	assert RAM(19620) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19620))))  severity failure;
	assert RAM(19621) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19621))))  severity failure;
	assert RAM(19622) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19622))))  severity failure;
	assert RAM(19623) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19623))))  severity failure;
	assert RAM(19624) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19624))))  severity failure;
	assert RAM(19625) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19625))))  severity failure;
	assert RAM(19626) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19626))))  severity failure;
	assert RAM(19627) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19627))))  severity failure;
	assert RAM(19628) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(19628))))  severity failure;
	assert RAM(19629) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19629))))  severity failure;
	assert RAM(19630) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19630))))  severity failure;
	assert RAM(19631) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19631))))  severity failure;
	assert RAM(19632) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19632))))  severity failure;
	assert RAM(19633) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19633))))  severity failure;
	assert RAM(19634) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19634))))  severity failure;
	assert RAM(19635) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19635))))  severity failure;
	assert RAM(19636) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19636))))  severity failure;
	assert RAM(19637) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19637))))  severity failure;
	assert RAM(19638) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19638))))  severity failure;
	assert RAM(19639) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19639))))  severity failure;
	assert RAM(19640) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19640))))  severity failure;
	assert RAM(19641) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19641))))  severity failure;
	assert RAM(19642) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(19642))))  severity failure;
	assert RAM(19643) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19643))))  severity failure;
	assert RAM(19644) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19644))))  severity failure;
	assert RAM(19645) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19645))))  severity failure;
	assert RAM(19646) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19646))))  severity failure;
	assert RAM(19647) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(19647))))  severity failure;
	assert RAM(19648) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19648))))  severity failure;
	assert RAM(19649) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(19649))))  severity failure;
	assert RAM(19650) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19650))))  severity failure;
	assert RAM(19651) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19651))))  severity failure;
	assert RAM(19652) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19652))))  severity failure;
	assert RAM(19653) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19653))))  severity failure;
	assert RAM(19654) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19654))))  severity failure;
	assert RAM(19655) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19655))))  severity failure;
	assert RAM(19656) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19656))))  severity failure;
	assert RAM(19657) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(19657))))  severity failure;
	assert RAM(19658) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19658))))  severity failure;
	assert RAM(19659) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19659))))  severity failure;
	assert RAM(19660) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19660))))  severity failure;
	assert RAM(19661) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19661))))  severity failure;
	assert RAM(19662) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19662))))  severity failure;
	assert RAM(19663) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19663))))  severity failure;
	assert RAM(19664) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19664))))  severity failure;
	assert RAM(19665) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19665))))  severity failure;
	assert RAM(19666) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(19666))))  severity failure;
	assert RAM(19667) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19667))))  severity failure;
	assert RAM(19668) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19668))))  severity failure;
	assert RAM(19669) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19669))))  severity failure;
	assert RAM(19670) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(19670))))  severity failure;
	assert RAM(19671) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19671))))  severity failure;
	assert RAM(19672) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19672))))  severity failure;
	assert RAM(19673) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19673))))  severity failure;
	assert RAM(19674) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19674))))  severity failure;
	assert RAM(19675) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19675))))  severity failure;
	assert RAM(19676) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19676))))  severity failure;
	assert RAM(19677) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19677))))  severity failure;
	assert RAM(19678) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(19678))))  severity failure;
	assert RAM(19679) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19679))))  severity failure;
	assert RAM(19680) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19680))))  severity failure;
	assert RAM(19681) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19681))))  severity failure;
	assert RAM(19682) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19682))))  severity failure;
	assert RAM(19683) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19683))))  severity failure;
	assert RAM(19684) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19684))))  severity failure;
	assert RAM(19685) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19685))))  severity failure;
	assert RAM(19686) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19686))))  severity failure;
	assert RAM(19687) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19687))))  severity failure;
	assert RAM(19688) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19688))))  severity failure;
	assert RAM(19689) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19689))))  severity failure;
	assert RAM(19690) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19690))))  severity failure;
	assert RAM(19691) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19691))))  severity failure;
	assert RAM(19692) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19692))))  severity failure;
	assert RAM(19693) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19693))))  severity failure;
	assert RAM(19694) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19694))))  severity failure;
	assert RAM(19695) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(19695))))  severity failure;
	assert RAM(19696) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19696))))  severity failure;
	assert RAM(19697) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19697))))  severity failure;
	assert RAM(19698) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19698))))  severity failure;
	assert RAM(19699) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(19699))))  severity failure;
	assert RAM(19700) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19700))))  severity failure;
	assert RAM(19701) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19701))))  severity failure;
	assert RAM(19702) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19702))))  severity failure;
	assert RAM(19703) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19703))))  severity failure;
	assert RAM(19704) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19704))))  severity failure;
	assert RAM(19705) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19705))))  severity failure;
	assert RAM(19706) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19706))))  severity failure;
	assert RAM(19707) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19707))))  severity failure;
	assert RAM(19708) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19708))))  severity failure;
	assert RAM(19709) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19709))))  severity failure;
	assert RAM(19710) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19710))))  severity failure;
	assert RAM(19711) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(19711))))  severity failure;
	assert RAM(19712) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19712))))  severity failure;
	assert RAM(19713) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19713))))  severity failure;
	assert RAM(19714) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19714))))  severity failure;
	assert RAM(19715) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19715))))  severity failure;
	assert RAM(19716) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(19716))))  severity failure;
	assert RAM(19717) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19717))))  severity failure;
	assert RAM(19718) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19718))))  severity failure;
	assert RAM(19719) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19719))))  severity failure;
	assert RAM(19720) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19720))))  severity failure;
	assert RAM(19721) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19721))))  severity failure;
	assert RAM(19722) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19722))))  severity failure;
	assert RAM(19723) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19723))))  severity failure;
	assert RAM(19724) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19724))))  severity failure;
	assert RAM(19725) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19725))))  severity failure;
	assert RAM(19726) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19726))))  severity failure;
	assert RAM(19727) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19727))))  severity failure;
	assert RAM(19728) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19728))))  severity failure;
	assert RAM(19729) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19729))))  severity failure;
	assert RAM(19730) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19730))))  severity failure;
	assert RAM(19731) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19731))))  severity failure;
	assert RAM(19732) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19732))))  severity failure;
	assert RAM(19733) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19733))))  severity failure;
	assert RAM(19734) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19734))))  severity failure;
	assert RAM(19735) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19735))))  severity failure;
	assert RAM(19736) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19736))))  severity failure;
	assert RAM(19737) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19737))))  severity failure;
	assert RAM(19738) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19738))))  severity failure;
	assert RAM(19739) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19739))))  severity failure;
	assert RAM(19740) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19740))))  severity failure;
	assert RAM(19741) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19741))))  severity failure;
	assert RAM(19742) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19742))))  severity failure;
	assert RAM(19743) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19743))))  severity failure;
	assert RAM(19744) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19744))))  severity failure;
	assert RAM(19745) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19745))))  severity failure;
	assert RAM(19746) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19746))))  severity failure;
	assert RAM(19747) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19747))))  severity failure;
	assert RAM(19748) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19748))))  severity failure;
	assert RAM(19749) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19749))))  severity failure;
	assert RAM(19750) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19750))))  severity failure;
	assert RAM(19751) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19751))))  severity failure;
	assert RAM(19752) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19752))))  severity failure;
	assert RAM(19753) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19753))))  severity failure;
	assert RAM(19754) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19754))))  severity failure;
	assert RAM(19755) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19755))))  severity failure;
	assert RAM(19756) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(19756))))  severity failure;
	assert RAM(19757) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(19757))))  severity failure;
	assert RAM(19758) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19758))))  severity failure;
	assert RAM(19759) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19759))))  severity failure;
	assert RAM(19760) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19760))))  severity failure;
	assert RAM(19761) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19761))))  severity failure;
	assert RAM(19762) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19762))))  severity failure;
	assert RAM(19763) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19763))))  severity failure;
	assert RAM(19764) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19764))))  severity failure;
	assert RAM(19765) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19765))))  severity failure;
	assert RAM(19766) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19766))))  severity failure;
	assert RAM(19767) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19767))))  severity failure;
	assert RAM(19768) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19768))))  severity failure;
	assert RAM(19769) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(19769))))  severity failure;
	assert RAM(19770) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(19770))))  severity failure;
	assert RAM(19771) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19771))))  severity failure;
	assert RAM(19772) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19772))))  severity failure;
	assert RAM(19773) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19773))))  severity failure;
	assert RAM(19774) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19774))))  severity failure;
	assert RAM(19775) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19775))))  severity failure;
	assert RAM(19776) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19776))))  severity failure;
	assert RAM(19777) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19777))))  severity failure;
	assert RAM(19778) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19778))))  severity failure;
	assert RAM(19779) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19779))))  severity failure;
	assert RAM(19780) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19780))))  severity failure;
	assert RAM(19781) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(19781))))  severity failure;
	assert RAM(19782) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19782))))  severity failure;
	assert RAM(19783) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19783))))  severity failure;
	assert RAM(19784) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19784))))  severity failure;
	assert RAM(19785) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19785))))  severity failure;
	assert RAM(19786) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19786))))  severity failure;
	assert RAM(19787) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19787))))  severity failure;
	assert RAM(19788) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19788))))  severity failure;
	assert RAM(19789) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19789))))  severity failure;
	assert RAM(19790) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(19790))))  severity failure;
	assert RAM(19791) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19791))))  severity failure;
	assert RAM(19792) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19792))))  severity failure;
	assert RAM(19793) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19793))))  severity failure;
	assert RAM(19794) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19794))))  severity failure;
	assert RAM(19795) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19795))))  severity failure;
	assert RAM(19796) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19796))))  severity failure;
	assert RAM(19797) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19797))))  severity failure;
	assert RAM(19798) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19798))))  severity failure;
	assert RAM(19799) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(19799))))  severity failure;
	assert RAM(19800) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19800))))  severity failure;
	assert RAM(19801) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19801))))  severity failure;
	assert RAM(19802) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19802))))  severity failure;
	assert RAM(19803) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19803))))  severity failure;
	assert RAM(19804) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19804))))  severity failure;
	assert RAM(19805) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19805))))  severity failure;
	assert RAM(19806) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19806))))  severity failure;
	assert RAM(19807) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19807))))  severity failure;
	assert RAM(19808) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(19808))))  severity failure;
	assert RAM(19809) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19809))))  severity failure;
	assert RAM(19810) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19810))))  severity failure;
	assert RAM(19811) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(19811))))  severity failure;
	assert RAM(19812) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19812))))  severity failure;
	assert RAM(19813) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19813))))  severity failure;
	assert RAM(19814) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19814))))  severity failure;
	assert RAM(19815) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(19815))))  severity failure;
	assert RAM(19816) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19816))))  severity failure;
	assert RAM(19817) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19817))))  severity failure;
	assert RAM(19818) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19818))))  severity failure;
	assert RAM(19819) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19819))))  severity failure;
	assert RAM(19820) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19820))))  severity failure;
	assert RAM(19821) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19821))))  severity failure;
	assert RAM(19822) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19822))))  severity failure;
	assert RAM(19823) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19823))))  severity failure;
	assert RAM(19824) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19824))))  severity failure;
	assert RAM(19825) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19825))))  severity failure;
	assert RAM(19826) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19826))))  severity failure;
	assert RAM(19827) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19827))))  severity failure;
	assert RAM(19828) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19828))))  severity failure;
	assert RAM(19829) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19829))))  severity failure;
	assert RAM(19830) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19830))))  severity failure;
	assert RAM(19831) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19831))))  severity failure;
	assert RAM(19832) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19832))))  severity failure;
	assert RAM(19833) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19833))))  severity failure;
	assert RAM(19834) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19834))))  severity failure;
	assert RAM(19835) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(19835))))  severity failure;
	assert RAM(19836) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19836))))  severity failure;
	assert RAM(19837) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19837))))  severity failure;
	assert RAM(19838) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(19838))))  severity failure;
	assert RAM(19839) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19839))))  severity failure;
	assert RAM(19840) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19840))))  severity failure;
	assert RAM(19841) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19841))))  severity failure;
	assert RAM(19842) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19842))))  severity failure;
	assert RAM(19843) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19843))))  severity failure;
	assert RAM(19844) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19844))))  severity failure;
	assert RAM(19845) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19845))))  severity failure;
	assert RAM(19846) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19846))))  severity failure;
	assert RAM(19847) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19847))))  severity failure;
	assert RAM(19848) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19848))))  severity failure;
	assert RAM(19849) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19849))))  severity failure;
	assert RAM(19850) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19850))))  severity failure;
	assert RAM(19851) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19851))))  severity failure;
	assert RAM(19852) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19852))))  severity failure;
	assert RAM(19853) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19853))))  severity failure;
	assert RAM(19854) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19854))))  severity failure;
	assert RAM(19855) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19855))))  severity failure;
	assert RAM(19856) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19856))))  severity failure;
	assert RAM(19857) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19857))))  severity failure;
	assert RAM(19858) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19858))))  severity failure;
	assert RAM(19859) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19859))))  severity failure;
	assert RAM(19860) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(19860))))  severity failure;
	assert RAM(19861) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19861))))  severity failure;
	assert RAM(19862) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19862))))  severity failure;
	assert RAM(19863) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19863))))  severity failure;
	assert RAM(19864) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19864))))  severity failure;
	assert RAM(19865) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19865))))  severity failure;
	assert RAM(19866) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(19866))))  severity failure;
	assert RAM(19867) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19867))))  severity failure;
	assert RAM(19868) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19868))))  severity failure;
	assert RAM(19869) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19869))))  severity failure;
	assert RAM(19870) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19870))))  severity failure;
	assert RAM(19871) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(19871))))  severity failure;
	assert RAM(19872) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19872))))  severity failure;
	assert RAM(19873) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19873))))  severity failure;
	assert RAM(19874) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19874))))  severity failure;
	assert RAM(19875) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19875))))  severity failure;
	assert RAM(19876) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19876))))  severity failure;
	assert RAM(19877) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19877))))  severity failure;
	assert RAM(19878) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19878))))  severity failure;
	assert RAM(19879) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19879))))  severity failure;
	assert RAM(19880) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(19880))))  severity failure;
	assert RAM(19881) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(19881))))  severity failure;
	assert RAM(19882) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19882))))  severity failure;
	assert RAM(19883) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(19883))))  severity failure;
	assert RAM(19884) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19884))))  severity failure;
	assert RAM(19885) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19885))))  severity failure;
	assert RAM(19886) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19886))))  severity failure;
	assert RAM(19887) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(19887))))  severity failure;
	assert RAM(19888) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19888))))  severity failure;
	assert RAM(19889) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19889))))  severity failure;
	assert RAM(19890) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19890))))  severity failure;
	assert RAM(19891) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19891))))  severity failure;
	assert RAM(19892) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19892))))  severity failure;
	assert RAM(19893) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19893))))  severity failure;
	assert RAM(19894) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19894))))  severity failure;
	assert RAM(19895) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19895))))  severity failure;
	assert RAM(19896) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19896))))  severity failure;
	assert RAM(19897) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(19897))))  severity failure;
	assert RAM(19898) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19898))))  severity failure;
	assert RAM(19899) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(19899))))  severity failure;
	assert RAM(19900) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19900))))  severity failure;
	assert RAM(19901) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19901))))  severity failure;
	assert RAM(19902) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19902))))  severity failure;
	assert RAM(19903) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19903))))  severity failure;
	assert RAM(19904) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19904))))  severity failure;
	assert RAM(19905) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(19905))))  severity failure;
	assert RAM(19906) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19906))))  severity failure;
	assert RAM(19907) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19907))))  severity failure;
	assert RAM(19908) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19908))))  severity failure;
	assert RAM(19909) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19909))))  severity failure;
	assert RAM(19910) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19910))))  severity failure;
	assert RAM(19911) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(19911))))  severity failure;
	assert RAM(19912) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19912))))  severity failure;
	assert RAM(19913) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19913))))  severity failure;
	assert RAM(19914) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19914))))  severity failure;
	assert RAM(19915) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19915))))  severity failure;
	assert RAM(19916) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19916))))  severity failure;
	assert RAM(19917) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(19917))))  severity failure;
	assert RAM(19918) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19918))))  severity failure;
	assert RAM(19919) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19919))))  severity failure;
	assert RAM(19920) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19920))))  severity failure;
	assert RAM(19921) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(19921))))  severity failure;
	assert RAM(19922) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19922))))  severity failure;
	assert RAM(19923) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19923))))  severity failure;
	assert RAM(19924) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19924))))  severity failure;
	assert RAM(19925) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19925))))  severity failure;
	assert RAM(19926) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19926))))  severity failure;
	assert RAM(19927) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19927))))  severity failure;
	assert RAM(19928) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19928))))  severity failure;
	assert RAM(19929) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19929))))  severity failure;
	assert RAM(19930) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19930))))  severity failure;
	assert RAM(19931) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19931))))  severity failure;
	assert RAM(19932) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19932))))  severity failure;
	assert RAM(19933) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19933))))  severity failure;
	assert RAM(19934) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19934))))  severity failure;
	assert RAM(19935) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19935))))  severity failure;
	assert RAM(19936) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19936))))  severity failure;
	assert RAM(19937) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19937))))  severity failure;
	assert RAM(19938) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19938))))  severity failure;
	assert RAM(19939) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19939))))  severity failure;
	assert RAM(19940) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19940))))  severity failure;
	assert RAM(19941) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19941))))  severity failure;
	assert RAM(19942) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19942))))  severity failure;
	assert RAM(19943) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(19943))))  severity failure;
	assert RAM(19944) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19944))))  severity failure;
	assert RAM(19945) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19945))))  severity failure;
	assert RAM(19946) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19946))))  severity failure;
	assert RAM(19947) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(19947))))  severity failure;
	assert RAM(19948) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19948))))  severity failure;
	assert RAM(19949) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19949))))  severity failure;
	assert RAM(19950) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19950))))  severity failure;
	assert RAM(19951) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19951))))  severity failure;
	assert RAM(19952) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19952))))  severity failure;
	assert RAM(19953) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19953))))  severity failure;
	assert RAM(19954) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19954))))  severity failure;
	assert RAM(19955) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19955))))  severity failure;
	assert RAM(19956) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19956))))  severity failure;
	assert RAM(19957) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19957))))  severity failure;
	assert RAM(19958) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(19958))))  severity failure;
	assert RAM(19959) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(19959))))  severity failure;
	assert RAM(19960) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19960))))  severity failure;
	assert RAM(19961) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19961))))  severity failure;
	assert RAM(19962) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(19962))))  severity failure;
	assert RAM(19963) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19963))))  severity failure;
	assert RAM(19964) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19964))))  severity failure;
	assert RAM(19965) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19965))))  severity failure;
	assert RAM(19966) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19966))))  severity failure;
	assert RAM(19967) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(19967))))  severity failure;
	assert RAM(19968) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19968))))  severity failure;
	assert RAM(19969) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19969))))  severity failure;
	assert RAM(19970) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19970))))  severity failure;
	assert RAM(19971) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19971))))  severity failure;
	assert RAM(19972) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19972))))  severity failure;
	assert RAM(19973) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19973))))  severity failure;
	assert RAM(19974) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19974))))  severity failure;
	assert RAM(19975) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19975))))  severity failure;
	assert RAM(19976) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19976))))  severity failure;
	assert RAM(19977) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19977))))  severity failure;
	assert RAM(19978) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19978))))  severity failure;
	assert RAM(19979) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19979))))  severity failure;
	assert RAM(19980) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19980))))  severity failure;
	assert RAM(19981) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19981))))  severity failure;
	assert RAM(19982) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19982))))  severity failure;
	assert RAM(19983) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19983))))  severity failure;
	assert RAM(19984) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19984))))  severity failure;
	assert RAM(19985) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19985))))  severity failure;
	assert RAM(19986) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19986))))  severity failure;
	assert RAM(19987) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19987))))  severity failure;
	assert RAM(19988) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19988))))  severity failure;
	assert RAM(19989) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19989))))  severity failure;
	assert RAM(19990) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19990))))  severity failure;
	assert RAM(19991) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19991))))  severity failure;
	assert RAM(19992) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19992))))  severity failure;
	assert RAM(19993) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19993))))  severity failure;
	assert RAM(19994) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19994))))  severity failure;
	assert RAM(19995) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19995))))  severity failure;
	assert RAM(19996) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19996))))  severity failure;
	assert RAM(19997) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19997))))  severity failure;
	assert RAM(19998) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19998))))  severity failure;
	assert RAM(19999) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19999))))  severity failure;
	assert RAM(20000) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20000))))  severity failure;
	assert RAM(20001) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20001))))  severity failure;
	assert RAM(20002) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20002))))  severity failure;
	assert RAM(20003) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20003))))  severity failure;
	assert RAM(20004) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(20004))))  severity failure;
	assert RAM(20005) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20005))))  severity failure;
	assert RAM(20006) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20006))))  severity failure;
	assert RAM(20007) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20007))))  severity failure;
	assert RAM(20008) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20008))))  severity failure;
	assert RAM(20009) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20009))))  severity failure;
	assert RAM(20010) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20010))))  severity failure;
	assert RAM(20011) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20011))))  severity failure;
	assert RAM(20012) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20012))))  severity failure;
	assert RAM(20013) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20013))))  severity failure;
	assert RAM(20014) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20014))))  severity failure;
	assert RAM(20015) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20015))))  severity failure;
	assert RAM(20016) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20016))))  severity failure;
	assert RAM(20017) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20017))))  severity failure;
	assert RAM(20018) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20018))))  severity failure;
	assert RAM(20019) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20019))))  severity failure;
	assert RAM(20020) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20020))))  severity failure;
	assert RAM(20021) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20021))))  severity failure;
	assert RAM(20022) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20022))))  severity failure;
	assert RAM(20023) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20023))))  severity failure;
	assert RAM(20024) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20024))))  severity failure;
	assert RAM(20025) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20025))))  severity failure;
	assert RAM(20026) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(20026))))  severity failure;
	assert RAM(20027) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20027))))  severity failure;
	assert RAM(20028) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20028))))  severity failure;
	assert RAM(20029) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20029))))  severity failure;
	assert RAM(20030) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20030))))  severity failure;
	assert RAM(20031) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20031))))  severity failure;
	assert RAM(20032) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20032))))  severity failure;
	assert RAM(20033) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20033))))  severity failure;
	assert RAM(20034) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20034))))  severity failure;
	assert RAM(20035) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20035))))  severity failure;
	assert RAM(20036) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20036))))  severity failure;
	assert RAM(20037) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20037))))  severity failure;
	assert RAM(20038) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20038))))  severity failure;
	assert RAM(20039) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20039))))  severity failure;
	assert RAM(20040) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20040))))  severity failure;
	assert RAM(20041) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20041))))  severity failure;
	assert RAM(20042) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20042))))  severity failure;
	assert RAM(20043) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20043))))  severity failure;
	assert RAM(20044) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20044))))  severity failure;
	assert RAM(20045) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20045))))  severity failure;
	assert RAM(20046) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(20046))))  severity failure;
	assert RAM(20047) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20047))))  severity failure;
	assert RAM(20048) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20048))))  severity failure;
	assert RAM(20049) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20049))))  severity failure;
	assert RAM(20050) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20050))))  severity failure;
	assert RAM(20051) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20051))))  severity failure;
	assert RAM(20052) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(20052))))  severity failure;
	assert RAM(20053) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20053))))  severity failure;
	assert RAM(20054) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20054))))  severity failure;
	assert RAM(20055) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20055))))  severity failure;
	assert RAM(20056) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20056))))  severity failure;
	assert RAM(20057) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20057))))  severity failure;
	assert RAM(20058) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20058))))  severity failure;
	assert RAM(20059) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20059))))  severity failure;
	assert RAM(20060) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20060))))  severity failure;
	assert RAM(20061) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20061))))  severity failure;
	assert RAM(20062) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20062))))  severity failure;
	assert RAM(20063) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20063))))  severity failure;
	assert RAM(20064) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20064))))  severity failure;
	assert RAM(20065) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20065))))  severity failure;
	assert RAM(20066) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(20066))))  severity failure;
	assert RAM(20067) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20067))))  severity failure;
	assert RAM(20068) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20068))))  severity failure;
	assert RAM(20069) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20069))))  severity failure;
	assert RAM(20070) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20070))))  severity failure;
	assert RAM(20071) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20071))))  severity failure;
	assert RAM(20072) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20072))))  severity failure;
	assert RAM(20073) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20073))))  severity failure;
	assert RAM(20074) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(20074))))  severity failure;
	assert RAM(20075) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20075))))  severity failure;
	assert RAM(20076) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20076))))  severity failure;
	assert RAM(20077) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20077))))  severity failure;
	assert RAM(20078) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20078))))  severity failure;
	assert RAM(20079) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20079))))  severity failure;
	assert RAM(20080) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20080))))  severity failure;
	assert RAM(20081) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(20081))))  severity failure;
	assert RAM(20082) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(20082))))  severity failure;
	assert RAM(20083) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20083))))  severity failure;
	assert RAM(20084) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20084))))  severity failure;
	assert RAM(20085) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20085))))  severity failure;
	assert RAM(20086) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20086))))  severity failure;
	assert RAM(20087) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20087))))  severity failure;
	assert RAM(20088) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20088))))  severity failure;
	assert RAM(20089) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20089))))  severity failure;
	assert RAM(20090) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20090))))  severity failure;
	assert RAM(20091) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20091))))  severity failure;
	assert RAM(20092) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(20092))))  severity failure;
	assert RAM(20093) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20093))))  severity failure;
	assert RAM(20094) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20094))))  severity failure;
	assert RAM(20095) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20095))))  severity failure;
	assert RAM(20096) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20096))))  severity failure;
	assert RAM(20097) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20097))))  severity failure;
	assert RAM(20098) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20098))))  severity failure;
	assert RAM(20099) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20099))))  severity failure;
	assert RAM(20100) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20100))))  severity failure;
	assert RAM(20101) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20101))))  severity failure;
	assert RAM(20102) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20102))))  severity failure;
	assert RAM(20103) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20103))))  severity failure;
	assert RAM(20104) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20104))))  severity failure;
	assert RAM(20105) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20105))))  severity failure;
	assert RAM(20106) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20106))))  severity failure;
	assert RAM(20107) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20107))))  severity failure;
	assert RAM(20108) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20108))))  severity failure;
	assert RAM(20109) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20109))))  severity failure;
	assert RAM(20110) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(20110))))  severity failure;
	assert RAM(20111) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20111))))  severity failure;
	assert RAM(20112) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20112))))  severity failure;
	assert RAM(20113) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20113))))  severity failure;
	assert RAM(20114) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20114))))  severity failure;
	assert RAM(20115) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20115))))  severity failure;
	assert RAM(20116) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20116))))  severity failure;
	assert RAM(20117) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20117))))  severity failure;
	assert RAM(20118) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20118))))  severity failure;
	assert RAM(20119) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20119))))  severity failure;
	assert RAM(20120) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(20120))))  severity failure;
	assert RAM(20121) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20121))))  severity failure;
	assert RAM(20122) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20122))))  severity failure;
	assert RAM(20123) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20123))))  severity failure;
	assert RAM(20124) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20124))))  severity failure;
	assert RAM(20125) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20125))))  severity failure;
	assert RAM(20126) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20126))))  severity failure;
	assert RAM(20127) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20127))))  severity failure;
	assert RAM(20128) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20128))))  severity failure;
	assert RAM(20129) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20129))))  severity failure;
	assert RAM(20130) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20130))))  severity failure;
	assert RAM(20131) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20131))))  severity failure;
	assert RAM(20132) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20132))))  severity failure;
	assert RAM(20133) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20133))))  severity failure;
	assert RAM(20134) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20134))))  severity failure;
	assert RAM(20135) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20135))))  severity failure;
	assert RAM(20136) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20136))))  severity failure;
	assert RAM(20137) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20137))))  severity failure;
	assert RAM(20138) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20138))))  severity failure;
	assert RAM(20139) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20139))))  severity failure;
	assert RAM(20140) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20140))))  severity failure;
	assert RAM(20141) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20141))))  severity failure;
	assert RAM(20142) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20142))))  severity failure;
	assert RAM(20143) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20143))))  severity failure;
	assert RAM(20144) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20144))))  severity failure;
	assert RAM(20145) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(20145))))  severity failure;
	assert RAM(20146) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20146))))  severity failure;
	assert RAM(20147) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20147))))  severity failure;
	assert RAM(20148) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20148))))  severity failure;
	assert RAM(20149) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20149))))  severity failure;
	assert RAM(20150) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20150))))  severity failure;
	assert RAM(20151) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20151))))  severity failure;
	assert RAM(20152) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20152))))  severity failure;
	assert RAM(20153) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20153))))  severity failure;
	assert RAM(20154) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20154))))  severity failure;
	assert RAM(20155) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20155))))  severity failure;
	assert RAM(20156) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20156))))  severity failure;
	assert RAM(20157) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20157))))  severity failure;
	assert RAM(20158) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20158))))  severity failure;
	assert RAM(20159) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20159))))  severity failure;
	assert RAM(20160) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20160))))  severity failure;
	assert RAM(20161) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20161))))  severity failure;
	assert RAM(20162) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20162))))  severity failure;
	assert RAM(20163) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20163))))  severity failure;
	assert RAM(20164) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20164))))  severity failure;
	assert RAM(20165) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20165))))  severity failure;
	assert RAM(20166) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20166))))  severity failure;
	assert RAM(20167) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20167))))  severity failure;
	assert RAM(20168) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20168))))  severity failure;
	assert RAM(20169) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20169))))  severity failure;
	assert RAM(20170) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20170))))  severity failure;
	assert RAM(20171) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20171))))  severity failure;
	assert RAM(20172) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20172))))  severity failure;
	assert RAM(20173) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20173))))  severity failure;
	assert RAM(20174) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20174))))  severity failure;
	assert RAM(20175) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20175))))  severity failure;
	assert RAM(20176) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20176))))  severity failure;
	assert RAM(20177) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20177))))  severity failure;
	assert RAM(20178) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(20178))))  severity failure;
	assert RAM(20179) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(20179))))  severity failure;
	assert RAM(20180) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20180))))  severity failure;
	assert RAM(20181) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20181))))  severity failure;
	assert RAM(20182) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20182))))  severity failure;
	assert RAM(20183) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20183))))  severity failure;
	assert RAM(20184) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(20184))))  severity failure;
	assert RAM(20185) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20185))))  severity failure;
	assert RAM(20186) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20186))))  severity failure;
	assert RAM(20187) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20187))))  severity failure;
	assert RAM(20188) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(20188))))  severity failure;
	assert RAM(20189) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(20189))))  severity failure;
	assert RAM(20190) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20190))))  severity failure;
	assert RAM(20191) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20191))))  severity failure;
	assert RAM(20192) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20192))))  severity failure;
	assert RAM(20193) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20193))))  severity failure;
	assert RAM(20194) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20194))))  severity failure;
	assert RAM(20195) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20195))))  severity failure;
	assert RAM(20196) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20196))))  severity failure;
	assert RAM(20197) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20197))))  severity failure;
	assert RAM(20198) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20198))))  severity failure;
	assert RAM(20199) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20199))))  severity failure;
	assert RAM(20200) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20200))))  severity failure;
	assert RAM(20201) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20201))))  severity failure;
	assert RAM(20202) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20202))))  severity failure;
	assert RAM(20203) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20203))))  severity failure;
	assert RAM(20204) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20204))))  severity failure;
	assert RAM(20205) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20205))))  severity failure;
	assert RAM(20206) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20206))))  severity failure;
	assert RAM(20207) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20207))))  severity failure;
	assert RAM(20208) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20208))))  severity failure;
	assert RAM(20209) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20209))))  severity failure;
	assert RAM(20210) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(20210))))  severity failure;
	assert RAM(20211) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(20211))))  severity failure;
	assert RAM(20212) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20212))))  severity failure;
	assert RAM(20213) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20213))))  severity failure;
	assert RAM(20214) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20214))))  severity failure;
	assert RAM(20215) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20215))))  severity failure;
	assert RAM(20216) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(20216))))  severity failure;
	assert RAM(20217) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20217))))  severity failure;
	assert RAM(20218) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20218))))  severity failure;
	assert RAM(20219) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20219))))  severity failure;
	assert RAM(20220) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(20220))))  severity failure;
	assert RAM(20221) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20221))))  severity failure;
	assert RAM(20222) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20222))))  severity failure;
	assert RAM(20223) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20223))))  severity failure;
	assert RAM(20224) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20224))))  severity failure;
	assert RAM(20225) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(20225))))  severity failure;
	assert RAM(20226) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20226))))  severity failure;
	assert RAM(20227) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20227))))  severity failure;
	assert RAM(20228) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(20228))))  severity failure;
	assert RAM(20229) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20229))))  severity failure;
	assert RAM(20230) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20230))))  severity failure;
	assert RAM(20231) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(20231))))  severity failure;
	assert RAM(20232) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20232))))  severity failure;
	assert RAM(20233) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20233))))  severity failure;
	assert RAM(20234) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20234))))  severity failure;
	assert RAM(20235) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20235))))  severity failure;
	assert RAM(20236) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20236))))  severity failure;
	assert RAM(20237) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20237))))  severity failure;
	assert RAM(20238) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20238))))  severity failure;
	assert RAM(20239) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20239))))  severity failure;
	assert RAM(20240) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20240))))  severity failure;
	assert RAM(20241) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20241))))  severity failure;
	assert RAM(20242) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(20242))))  severity failure;
	assert RAM(20243) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20243))))  severity failure;
	assert RAM(20244) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20244))))  severity failure;
	assert RAM(20245) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20245))))  severity failure;
	assert RAM(20246) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20246))))  severity failure;
	assert RAM(20247) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20247))))  severity failure;
	assert RAM(20248) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20248))))  severity failure;
	assert RAM(20249) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20249))))  severity failure;
	assert RAM(20250) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20250))))  severity failure;
	assert RAM(20251) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20251))))  severity failure;
	assert RAM(20252) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20252))))  severity failure;
	assert RAM(20253) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(20253))))  severity failure;
	assert RAM(20254) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20254))))  severity failure;
	assert RAM(20255) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20255))))  severity failure;
	assert RAM(20256) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(20256))))  severity failure;
	assert RAM(20257) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20257))))  severity failure;
	assert RAM(20258) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20258))))  severity failure;
	assert RAM(20259) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20259))))  severity failure;
	assert RAM(20260) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20260))))  severity failure;
	assert RAM(20261) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20261))))  severity failure;
	assert RAM(20262) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20262))))  severity failure;
	assert RAM(20263) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20263))))  severity failure;
	assert RAM(20264) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20264))))  severity failure;
	assert RAM(20265) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20265))))  severity failure;
	assert RAM(20266) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20266))))  severity failure;
	assert RAM(20267) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(20267))))  severity failure;
	assert RAM(20268) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20268))))  severity failure;
	assert RAM(20269) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20269))))  severity failure;
	assert RAM(20270) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20270))))  severity failure;
	assert RAM(20271) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20271))))  severity failure;
	assert RAM(20272) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20272))))  severity failure;
	assert RAM(20273) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20273))))  severity failure;
	assert RAM(20274) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20274))))  severity failure;
	assert RAM(20275) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20275))))  severity failure;
	assert RAM(20276) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20276))))  severity failure;
	assert RAM(20277) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(20277))))  severity failure;
	assert RAM(20278) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20278))))  severity failure;
	assert RAM(20279) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20279))))  severity failure;
	assert RAM(20280) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20280))))  severity failure;
	assert RAM(20281) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20281))))  severity failure;
	assert RAM(20282) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20282))))  severity failure;
	assert RAM(20283) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(20283))))  severity failure;
	assert RAM(20284) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20284))))  severity failure;
	assert RAM(20285) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20285))))  severity failure;
	assert RAM(20286) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20286))))  severity failure;
	assert RAM(20287) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20287))))  severity failure;
	assert RAM(20288) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(20288))))  severity failure;
	assert RAM(20289) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20289))))  severity failure;
	assert RAM(20290) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20290))))  severity failure;
	assert RAM(20291) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20291))))  severity failure;
	assert RAM(20292) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20292))))  severity failure;
	assert RAM(20293) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20293))))  severity failure;
	assert RAM(20294) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20294))))  severity failure;
	assert RAM(20295) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20295))))  severity failure;
	assert RAM(20296) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20296))))  severity failure;
	assert RAM(20297) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20297))))  severity failure;
	assert RAM(20298) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20298))))  severity failure;
	assert RAM(20299) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20299))))  severity failure;
	assert RAM(20300) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(20300))))  severity failure;
	assert RAM(20301) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20301))))  severity failure;
	assert RAM(20302) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20302))))  severity failure;
	assert RAM(20303) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20303))))  severity failure;
	assert RAM(20304) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20304))))  severity failure;
	assert RAM(20305) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20305))))  severity failure;
	assert RAM(20306) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20306))))  severity failure;
	assert RAM(20307) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20307))))  severity failure;
	assert RAM(20308) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20308))))  severity failure;
	assert RAM(20309) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(20309))))  severity failure;
	assert RAM(20310) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20310))))  severity failure;
	assert RAM(20311) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20311))))  severity failure;
	assert RAM(20312) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20312))))  severity failure;
	assert RAM(20313) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20313))))  severity failure;
	assert RAM(20314) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20314))))  severity failure;
	assert RAM(20315) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20315))))  severity failure;
	assert RAM(20316) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(20316))))  severity failure;
	assert RAM(20317) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20317))))  severity failure;
	assert RAM(20318) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(20318))))  severity failure;
	assert RAM(20319) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20319))))  severity failure;
	assert RAM(20320) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20320))))  severity failure;
	assert RAM(20321) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20321))))  severity failure;
	assert RAM(20322) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20322))))  severity failure;
	assert RAM(20323) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(20323))))  severity failure;
	assert RAM(20324) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20324))))  severity failure;
	assert RAM(20325) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20325))))  severity failure;
	assert RAM(20326) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20326))))  severity failure;
	assert RAM(20327) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20327))))  severity failure;
	assert RAM(20328) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20328))))  severity failure;
	assert RAM(20329) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20329))))  severity failure;
	assert RAM(20330) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20330))))  severity failure;
	assert RAM(20331) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20331))))  severity failure;
	assert RAM(20332) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20332))))  severity failure;
	assert RAM(20333) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20333))))  severity failure;
	assert RAM(20334) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(20334))))  severity failure;
	assert RAM(20335) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20335))))  severity failure;
	assert RAM(20336) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20336))))  severity failure;
	assert RAM(20337) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20337))))  severity failure;
	assert RAM(20338) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20338))))  severity failure;
	assert RAM(20339) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(20339))))  severity failure;
	assert RAM(20340) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20340))))  severity failure;
	assert RAM(20341) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20341))))  severity failure;
	assert RAM(20342) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20342))))  severity failure;
	assert RAM(20343) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20343))))  severity failure;
	assert RAM(20344) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20344))))  severity failure;
	assert RAM(20345) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20345))))  severity failure;
	assert RAM(20346) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20346))))  severity failure;
	assert RAM(20347) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(20347))))  severity failure;
	assert RAM(20348) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20348))))  severity failure;
	assert RAM(20349) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20349))))  severity failure;
	assert RAM(20350) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20350))))  severity failure;
	assert RAM(20351) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(20351))))  severity failure;
	assert RAM(20352) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(20352))))  severity failure;
	assert RAM(20353) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20353))))  severity failure;
	assert RAM(20354) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20354))))  severity failure;
	assert RAM(20355) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20355))))  severity failure;
	assert RAM(20356) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(20356))))  severity failure;
	assert RAM(20357) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20357))))  severity failure;
	assert RAM(20358) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20358))))  severity failure;
	assert RAM(20359) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20359))))  severity failure;
	assert RAM(20360) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20360))))  severity failure;
	assert RAM(20361) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20361))))  severity failure;
	assert RAM(20362) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20362))))  severity failure;
	assert RAM(20363) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20363))))  severity failure;
	assert RAM(20364) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20364))))  severity failure;
	assert RAM(20365) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20365))))  severity failure;
	assert RAM(20366) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20366))))  severity failure;
	assert RAM(20367) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20367))))  severity failure;
	assert RAM(20368) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20368))))  severity failure;
	assert RAM(20369) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20369))))  severity failure;
	assert RAM(20370) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(20370))))  severity failure;
	assert RAM(20371) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20371))))  severity failure;
	assert RAM(20372) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20372))))  severity failure;
	assert RAM(20373) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20373))))  severity failure;
	assert RAM(20374) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20374))))  severity failure;
	assert RAM(20375) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(20375))))  severity failure;
	assert RAM(20376) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(20376))))  severity failure;
	assert RAM(20377) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20377))))  severity failure;
	assert RAM(20378) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20378))))  severity failure;
	assert RAM(20379) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20379))))  severity failure;
	assert RAM(20380) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20380))))  severity failure;
	assert RAM(20381) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20381))))  severity failure;
	assert RAM(20382) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20382))))  severity failure;
	assert RAM(20383) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20383))))  severity failure;
	assert RAM(20384) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(20384))))  severity failure;
	assert RAM(20385) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20385))))  severity failure;
	assert RAM(20386) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20386))))  severity failure;
	assert RAM(20387) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(20387))))  severity failure;
	assert RAM(20388) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20388))))  severity failure;
	assert RAM(20389) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(20389))))  severity failure;
	assert RAM(20390) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20390))))  severity failure;
	assert RAM(20391) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20391))))  severity failure;
	assert RAM(20392) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20392))))  severity failure;
	assert RAM(20393) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20393))))  severity failure;
	assert RAM(20394) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20394))))  severity failure;
	assert RAM(20395) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20395))))  severity failure;
	assert RAM(20396) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20396))))  severity failure;
	assert RAM(20397) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20397))))  severity failure;
	assert RAM(20398) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20398))))  severity failure;
	assert RAM(20399) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20399))))  severity failure;
	assert RAM(20400) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20400))))  severity failure;
	assert RAM(20401) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20401))))  severity failure;
	assert RAM(20402) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(20402))))  severity failure;
	assert RAM(20403) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20403))))  severity failure;
	assert RAM(20404) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20404))))  severity failure;
	assert RAM(20405) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20405))))  severity failure;
	assert RAM(20406) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20406))))  severity failure;
	assert RAM(20407) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20407))))  severity failure;
	assert RAM(20408) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20408))))  severity failure;
	assert RAM(20409) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20409))))  severity failure;
	assert RAM(20410) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(20410))))  severity failure;
	assert RAM(20411) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20411))))  severity failure;
	assert RAM(20412) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20412))))  severity failure;
	assert RAM(20413) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20413))))  severity failure;
	assert RAM(20414) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20414))))  severity failure;
	assert RAM(20415) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20415))))  severity failure;
	assert RAM(20416) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20416))))  severity failure;
	assert RAM(20417) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20417))))  severity failure;
	assert RAM(20418) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20418))))  severity failure;
	assert RAM(20419) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20419))))  severity failure;
	assert RAM(20420) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20420))))  severity failure;
	assert RAM(20421) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20421))))  severity failure;
	assert RAM(20422) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(20422))))  severity failure;
	assert RAM(20423) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20423))))  severity failure;
	assert RAM(20424) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20424))))  severity failure;
	assert RAM(20425) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20425))))  severity failure;
	assert RAM(20426) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20426))))  severity failure;
	assert RAM(20427) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20427))))  severity failure;
	assert RAM(20428) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20428))))  severity failure;
	assert RAM(20429) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20429))))  severity failure;
	assert RAM(20430) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20430))))  severity failure;
	assert RAM(20431) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20431))))  severity failure;
	assert RAM(20432) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20432))))  severity failure;
	assert RAM(20433) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20433))))  severity failure;
	assert RAM(20434) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(20434))))  severity failure;
	assert RAM(20435) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20435))))  severity failure;
	assert RAM(20436) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20436))))  severity failure;
	assert RAM(20437) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20437))))  severity failure;
	assert RAM(20438) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(20438))))  severity failure;
	assert RAM(20439) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20439))))  severity failure;
	assert RAM(20440) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20440))))  severity failure;
	assert RAM(20441) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20441))))  severity failure;
	assert RAM(20442) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(20442))))  severity failure;
	assert RAM(20443) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20443))))  severity failure;
	assert RAM(20444) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(20444))))  severity failure;
	assert RAM(20445) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20445))))  severity failure;
	assert RAM(20446) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20446))))  severity failure;
	assert RAM(20447) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20447))))  severity failure;
	assert RAM(20448) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20448))))  severity failure;
	assert RAM(20449) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20449))))  severity failure;
	assert RAM(20450) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20450))))  severity failure;
	assert RAM(20451) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20451))))  severity failure;
	assert RAM(20452) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(20452))))  severity failure;
	assert RAM(20453) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20453))))  severity failure;
	assert RAM(20454) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20454))))  severity failure;
	assert RAM(20455) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20455))))  severity failure;
	assert RAM(20456) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20456))))  severity failure;
	assert RAM(20457) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20457))))  severity failure;
	assert RAM(20458) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20458))))  severity failure;
	assert RAM(20459) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20459))))  severity failure;
	assert RAM(20460) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20460))))  severity failure;
	assert RAM(20461) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20461))))  severity failure;
	assert RAM(20462) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20462))))  severity failure;
	assert RAM(20463) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20463))))  severity failure;
	assert RAM(20464) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20464))))  severity failure;
	assert RAM(20465) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20465))))  severity failure;
	assert RAM(20466) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20466))))  severity failure;
	assert RAM(20467) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20467))))  severity failure;
	assert RAM(20468) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20468))))  severity failure;
	assert RAM(20469) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(20469))))  severity failure;
	assert RAM(20470) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(20470))))  severity failure;
	assert RAM(20471) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20471))))  severity failure;
	assert RAM(20472) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20472))))  severity failure;
	assert RAM(20473) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(20473))))  severity failure;
	assert RAM(20474) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20474))))  severity failure;
	assert RAM(20475) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20475))))  severity failure;
	assert RAM(20476) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20476))))  severity failure;
	assert RAM(20477) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20477))))  severity failure;
	assert RAM(20478) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20478))))  severity failure;
	assert RAM(20479) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20479))))  severity failure;
	assert RAM(20480) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20480))))  severity failure;
	assert RAM(20481) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20481))))  severity failure;
	assert RAM(20482) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20482))))  severity failure;
	assert RAM(20483) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20483))))  severity failure;
	assert RAM(20484) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20484))))  severity failure;
	assert RAM(20485) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20485))))  severity failure;
	assert RAM(20486) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20486))))  severity failure;
	assert RAM(20487) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20487))))  severity failure;
	assert RAM(20488) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(20488))))  severity failure;
	assert RAM(20489) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20489))))  severity failure;
	assert RAM(20490) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20490))))  severity failure;
	assert RAM(20491) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(20491))))  severity failure;
	assert RAM(20492) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20492))))  severity failure;
	assert RAM(20493) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20493))))  severity failure;
	assert RAM(20494) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20494))))  severity failure;
	assert RAM(20495) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20495))))  severity failure;
	assert RAM(20496) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20496))))  severity failure;
	assert RAM(20497) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20497))))  severity failure;
	assert RAM(20498) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20498))))  severity failure;
	assert RAM(20499) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20499))))  severity failure;
	assert RAM(20500) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20500))))  severity failure;
	assert RAM(20501) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20501))))  severity failure;
	assert RAM(20502) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20502))))  severity failure;
	assert RAM(20503) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20503))))  severity failure;
	assert RAM(20504) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20504))))  severity failure;
	assert RAM(20505) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20505))))  severity failure;
	assert RAM(20506) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20506))))  severity failure;
	assert RAM(20507) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20507))))  severity failure;
	assert RAM(20508) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20508))))  severity failure;
	assert RAM(20509) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20509))))  severity failure;
	assert RAM(20510) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20510))))  severity failure;
	assert RAM(20511) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20511))))  severity failure;
	assert RAM(20512) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(20512))))  severity failure;
	assert RAM(20513) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20513))))  severity failure;
	assert RAM(20514) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20514))))  severity failure;
	assert RAM(20515) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20515))))  severity failure;
	assert RAM(20516) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(20516))))  severity failure;
	assert RAM(20517) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20517))))  severity failure;
	assert RAM(20518) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20518))))  severity failure;
	assert RAM(20519) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(20519))))  severity failure;
	assert RAM(20520) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20520))))  severity failure;
	assert RAM(20521) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20521))))  severity failure;
	assert RAM(20522) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20522))))  severity failure;
	assert RAM(20523) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20523))))  severity failure;
	assert RAM(20524) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20524))))  severity failure;
	assert RAM(20525) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20525))))  severity failure;
	assert RAM(20526) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20526))))  severity failure;
	assert RAM(20527) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20527))))  severity failure;
	assert RAM(20528) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(20528))))  severity failure;
	assert RAM(20529) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20529))))  severity failure;
	assert RAM(20530) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20530))))  severity failure;
	assert RAM(20531) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20531))))  severity failure;
	assert RAM(20532) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20532))))  severity failure;
	assert RAM(20533) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20533))))  severity failure;
	assert RAM(20534) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20534))))  severity failure;
	assert RAM(20535) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20535))))  severity failure;
	assert RAM(20536) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20536))))  severity failure;
	assert RAM(20537) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20537))))  severity failure;
	assert RAM(20538) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20538))))  severity failure;
	assert RAM(20539) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(20539))))  severity failure;
	assert RAM(20540) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20540))))  severity failure;
	assert RAM(20541) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20541))))  severity failure;
	assert RAM(20542) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20542))))  severity failure;
	assert RAM(20543) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20543))))  severity failure;
	assert RAM(20544) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20544))))  severity failure;
	assert RAM(20545) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(20545))))  severity failure;
	assert RAM(20546) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20546))))  severity failure;
	assert RAM(20547) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20547))))  severity failure;
	assert RAM(20548) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20548))))  severity failure;
	assert RAM(20549) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20549))))  severity failure;
	assert RAM(20550) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20550))))  severity failure;
	assert RAM(20551) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20551))))  severity failure;
	assert RAM(20552) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20552))))  severity failure;
	assert RAM(20553) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20553))))  severity failure;
	assert RAM(20554) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20554))))  severity failure;
	assert RAM(20555) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20555))))  severity failure;
	assert RAM(20556) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20556))))  severity failure;
	assert RAM(20557) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(20557))))  severity failure;
	assert RAM(20558) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20558))))  severity failure;
	assert RAM(20559) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20559))))  severity failure;
	assert RAM(20560) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20560))))  severity failure;
	assert RAM(20561) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20561))))  severity failure;
	assert RAM(20562) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(20562))))  severity failure;
	assert RAM(20563) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(20563))))  severity failure;
	assert RAM(20564) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20564))))  severity failure;
	assert RAM(20565) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20565))))  severity failure;
	assert RAM(20566) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20566))))  severity failure;
	assert RAM(20567) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20567))))  severity failure;
	assert RAM(20568) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20568))))  severity failure;
	assert RAM(20569) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20569))))  severity failure;
	assert RAM(20570) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(20570))))  severity failure;
	assert RAM(20571) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20571))))  severity failure;
	assert RAM(20572) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20572))))  severity failure;
	assert RAM(20573) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(20573))))  severity failure;
	assert RAM(20574) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20574))))  severity failure;
	assert RAM(20575) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20575))))  severity failure;
	assert RAM(20576) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20576))))  severity failure;
	assert RAM(20577) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20577))))  severity failure;
	assert RAM(20578) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20578))))  severity failure;
	assert RAM(20579) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20579))))  severity failure;
	assert RAM(20580) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20580))))  severity failure;
	assert RAM(20581) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20581))))  severity failure;
	assert RAM(20582) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20582))))  severity failure;
	assert RAM(20583) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20583))))  severity failure;
	assert RAM(20584) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20584))))  severity failure;
	assert RAM(20585) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(20585))))  severity failure;
	assert RAM(20586) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20586))))  severity failure;
	assert RAM(20587) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(20587))))  severity failure;
	assert RAM(20588) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20588))))  severity failure;
	assert RAM(20589) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20589))))  severity failure;
	assert RAM(20590) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20590))))  severity failure;
	assert RAM(20591) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20591))))  severity failure;
	assert RAM(20592) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20592))))  severity failure;
	assert RAM(20593) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20593))))  severity failure;
	assert RAM(20594) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20594))))  severity failure;
	assert RAM(20595) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20595))))  severity failure;
	assert RAM(20596) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(20596))))  severity failure;
	assert RAM(20597) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20597))))  severity failure;
	assert RAM(20598) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20598))))  severity failure;
	assert RAM(20599) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(20599))))  severity failure;
	assert RAM(20600) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20600))))  severity failure;
	assert RAM(20601) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20601))))  severity failure;
	assert RAM(20602) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20602))))  severity failure;
	assert RAM(20603) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20603))))  severity failure;
	assert RAM(20604) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20604))))  severity failure;
	assert RAM(20605) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20605))))  severity failure;
	assert RAM(20606) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(20606))))  severity failure;
	assert RAM(20607) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20607))))  severity failure;
	assert RAM(20608) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20608))))  severity failure;
	assert RAM(20609) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20609))))  severity failure;
	assert RAM(20610) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20610))))  severity failure;
	assert RAM(20611) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20611))))  severity failure;
	assert RAM(20612) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20612))))  severity failure;
	assert RAM(20613) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20613))))  severity failure;
	assert RAM(20614) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20614))))  severity failure;
	assert RAM(20615) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20615))))  severity failure;
	assert RAM(20616) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20616))))  severity failure;
	assert RAM(20617) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(20617))))  severity failure;
	assert RAM(20618) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20618))))  severity failure;
	assert RAM(20619) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20619))))  severity failure;
	assert RAM(20620) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20620))))  severity failure;
	assert RAM(20621) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20621))))  severity failure;
	assert RAM(20622) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20622))))  severity failure;
	assert RAM(20623) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20623))))  severity failure;
	assert RAM(20624) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(20624))))  severity failure;
	assert RAM(20625) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(20625))))  severity failure;
	assert RAM(20626) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20626))))  severity failure;
	assert RAM(20627) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20627))))  severity failure;
	assert RAM(20628) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20628))))  severity failure;
	assert RAM(20629) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20629))))  severity failure;
	assert RAM(20630) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20630))))  severity failure;
	assert RAM(20631) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20631))))  severity failure;
	assert RAM(20632) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20632))))  severity failure;
	assert RAM(20633) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20633))))  severity failure;
	assert RAM(20634) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20634))))  severity failure;
	assert RAM(20635) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20635))))  severity failure;
	assert RAM(20636) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20636))))  severity failure;
	assert RAM(20637) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20637))))  severity failure;
	assert RAM(20638) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20638))))  severity failure;
	assert RAM(20639) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20639))))  severity failure;
	assert RAM(20640) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20640))))  severity failure;
	assert RAM(20641) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20641))))  severity failure;
	assert RAM(20642) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20642))))  severity failure;
	assert RAM(20643) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20643))))  severity failure;
	assert RAM(20644) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20644))))  severity failure;
	assert RAM(20645) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20645))))  severity failure;
	assert RAM(20646) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20646))))  severity failure;
	assert RAM(20647) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20647))))  severity failure;
	assert RAM(20648) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20648))))  severity failure;
	assert RAM(20649) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20649))))  severity failure;
	assert RAM(20650) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20650))))  severity failure;
	assert RAM(20651) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20651))))  severity failure;
	assert RAM(20652) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20652))))  severity failure;
	assert RAM(20653) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20653))))  severity failure;
	assert RAM(20654) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20654))))  severity failure;
	assert RAM(20655) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20655))))  severity failure;
	assert RAM(20656) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20656))))  severity failure;
	assert RAM(20657) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20657))))  severity failure;
	assert RAM(20658) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20658))))  severity failure;
	assert RAM(20659) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20659))))  severity failure;
	assert RAM(20660) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20660))))  severity failure;
	assert RAM(20661) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20661))))  severity failure;
	assert RAM(20662) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20662))))  severity failure;
	assert RAM(20663) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(20663))))  severity failure;
	assert RAM(20664) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20664))))  severity failure;
	assert RAM(20665) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20665))))  severity failure;
	assert RAM(20666) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20666))))  severity failure;
	assert RAM(20667) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20667))))  severity failure;
	assert RAM(20668) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20668))))  severity failure;
	assert RAM(20669) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20669))))  severity failure;
	assert RAM(20670) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20670))))  severity failure;
	assert RAM(20671) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20671))))  severity failure;
	assert RAM(20672) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20672))))  severity failure;
	assert RAM(20673) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20673))))  severity failure;
	assert RAM(20674) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(20674))))  severity failure;
	assert RAM(20675) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20675))))  severity failure;
	assert RAM(20676) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20676))))  severity failure;
	assert RAM(20677) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20677))))  severity failure;
	assert RAM(20678) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20678))))  severity failure;
	assert RAM(20679) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20679))))  severity failure;
	assert RAM(20680) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20680))))  severity failure;
	assert RAM(20681) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20681))))  severity failure;
	assert RAM(20682) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20682))))  severity failure;
	assert RAM(20683) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20683))))  severity failure;
	assert RAM(20684) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20684))))  severity failure;
	assert RAM(20685) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20685))))  severity failure;
	assert RAM(20686) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20686))))  severity failure;
	assert RAM(20687) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20687))))  severity failure;
	assert RAM(20688) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20688))))  severity failure;
	assert RAM(20689) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20689))))  severity failure;
	assert RAM(20690) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20690))))  severity failure;
	assert RAM(20691) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(20691))))  severity failure;
	assert RAM(20692) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20692))))  severity failure;
	assert RAM(20693) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20693))))  severity failure;
	assert RAM(20694) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20694))))  severity failure;
	assert RAM(20695) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20695))))  severity failure;
	assert RAM(20696) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20696))))  severity failure;
	assert RAM(20697) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20697))))  severity failure;
	assert RAM(20698) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20698))))  severity failure;
	assert RAM(20699) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20699))))  severity failure;
	assert RAM(20700) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20700))))  severity failure;
	assert RAM(20701) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20701))))  severity failure;
	assert RAM(20702) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20702))))  severity failure;
	assert RAM(20703) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20703))))  severity failure;
	assert RAM(20704) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20704))))  severity failure;
	assert RAM(20705) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20705))))  severity failure;
	assert RAM(20706) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20706))))  severity failure;
	assert RAM(20707) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20707))))  severity failure;
	assert RAM(20708) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20708))))  severity failure;
	assert RAM(20709) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20709))))  severity failure;
	assert RAM(20710) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20710))))  severity failure;
	assert RAM(20711) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20711))))  severity failure;
	assert RAM(20712) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20712))))  severity failure;
	assert RAM(20713) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20713))))  severity failure;
	assert RAM(20714) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20714))))  severity failure;
	assert RAM(20715) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20715))))  severity failure;
	assert RAM(20716) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20716))))  severity failure;
	assert RAM(20717) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20717))))  severity failure;
	assert RAM(20718) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(20718))))  severity failure;
	assert RAM(20719) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20719))))  severity failure;
	assert RAM(20720) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20720))))  severity failure;
	assert RAM(20721) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20721))))  severity failure;
	assert RAM(20722) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20722))))  severity failure;
	assert RAM(20723) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20723))))  severity failure;
	assert RAM(20724) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20724))))  severity failure;
	assert RAM(20725) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(20725))))  severity failure;
	assert RAM(20726) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20726))))  severity failure;
	assert RAM(20727) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20727))))  severity failure;
	assert RAM(20728) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20728))))  severity failure;
	assert RAM(20729) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20729))))  severity failure;
	assert RAM(20730) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20730))))  severity failure;
	assert RAM(20731) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20731))))  severity failure;
	assert RAM(20732) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20732))))  severity failure;
	assert RAM(20733) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20733))))  severity failure;
	assert RAM(20734) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20734))))  severity failure;
	assert RAM(20735) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20735))))  severity failure;
	assert RAM(20736) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20736))))  severity failure;
	assert RAM(20737) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20737))))  severity failure;
	assert RAM(20738) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(20738))))  severity failure;
	assert RAM(20739) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20739))))  severity failure;
	assert RAM(20740) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20740))))  severity failure;
	assert RAM(20741) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20741))))  severity failure;
	assert RAM(20742) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20742))))  severity failure;
	assert RAM(20743) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(20743))))  severity failure;
	assert RAM(20744) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20744))))  severity failure;
	assert RAM(20745) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20745))))  severity failure;
	assert RAM(20746) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20746))))  severity failure;
	assert RAM(20747) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20747))))  severity failure;
	assert RAM(20748) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20748))))  severity failure;
	assert RAM(20749) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20749))))  severity failure;
	assert RAM(20750) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20750))))  severity failure;
	assert RAM(20751) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20751))))  severity failure;
	assert RAM(20752) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(20752))))  severity failure;
	assert RAM(20753) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20753))))  severity failure;
	assert RAM(20754) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20754))))  severity failure;
	assert RAM(20755) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20755))))  severity failure;
	assert RAM(20756) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20756))))  severity failure;
	assert RAM(20757) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20757))))  severity failure;
	assert RAM(20758) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20758))))  severity failure;
	assert RAM(20759) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(20759))))  severity failure;
	assert RAM(20760) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(20760))))  severity failure;
	assert RAM(20761) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20761))))  severity failure;
	assert RAM(20762) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20762))))  severity failure;
	assert RAM(20763) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20763))))  severity failure;
	assert RAM(20764) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20764))))  severity failure;
	assert RAM(20765) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(20765))))  severity failure;
	assert RAM(20766) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20766))))  severity failure;
	assert RAM(20767) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(20767))))  severity failure;
	assert RAM(20768) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20768))))  severity failure;
	assert RAM(20769) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20769))))  severity failure;
	assert RAM(20770) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20770))))  severity failure;
	assert RAM(20771) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20771))))  severity failure;
	assert RAM(20772) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20772))))  severity failure;
	assert RAM(20773) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20773))))  severity failure;
	assert RAM(20774) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(20774))))  severity failure;
	assert RAM(20775) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20775))))  severity failure;
	assert RAM(20776) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20776))))  severity failure;
	assert RAM(20777) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20777))))  severity failure;
	assert RAM(20778) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20778))))  severity failure;
	assert RAM(20779) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20779))))  severity failure;
	assert RAM(20780) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20780))))  severity failure;
	assert RAM(20781) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20781))))  severity failure;
	assert RAM(20782) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20782))))  severity failure;
	assert RAM(20783) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20783))))  severity failure;
	assert RAM(20784) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20784))))  severity failure;
	assert RAM(20785) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20785))))  severity failure;
	assert RAM(20786) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20786))))  severity failure;
	assert RAM(20787) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20787))))  severity failure;
	assert RAM(20788) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20788))))  severity failure;
	assert RAM(20789) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20789))))  severity failure;
	assert RAM(20790) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20790))))  severity failure;
	assert RAM(20791) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(20791))))  severity failure;
	assert RAM(20792) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20792))))  severity failure;
	assert RAM(20793) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20793))))  severity failure;
	assert RAM(20794) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20794))))  severity failure;
	assert RAM(20795) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20795))))  severity failure;
	assert RAM(20796) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20796))))  severity failure;
	assert RAM(20797) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20797))))  severity failure;
	assert RAM(20798) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20798))))  severity failure;
	assert RAM(20799) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20799))))  severity failure;
	assert RAM(20800) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20800))))  severity failure;
	assert RAM(20801) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20801))))  severity failure;
	assert RAM(20802) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20802))))  severity failure;
	assert RAM(20803) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(20803))))  severity failure;
	assert RAM(20804) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20804))))  severity failure;
	assert RAM(20805) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20805))))  severity failure;
	assert RAM(20806) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20806))))  severity failure;
	assert RAM(20807) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20807))))  severity failure;
	assert RAM(20808) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20808))))  severity failure;
	assert RAM(20809) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20809))))  severity failure;
	assert RAM(20810) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20810))))  severity failure;
	assert RAM(20811) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20811))))  severity failure;
	assert RAM(20812) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20812))))  severity failure;
	assert RAM(20813) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20813))))  severity failure;
	assert RAM(20814) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20814))))  severity failure;
	assert RAM(20815) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20815))))  severity failure;
	assert RAM(20816) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20816))))  severity failure;
	assert RAM(20817) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20817))))  severity failure;
	assert RAM(20818) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20818))))  severity failure;
	assert RAM(20819) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20819))))  severity failure;
	assert RAM(20820) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20820))))  severity failure;
	assert RAM(20821) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(20821))))  severity failure;
	assert RAM(20822) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20822))))  severity failure;
	assert RAM(20823) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(20823))))  severity failure;
	assert RAM(20824) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20824))))  severity failure;
	assert RAM(20825) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20825))))  severity failure;
	assert RAM(20826) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20826))))  severity failure;
	assert RAM(20827) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20827))))  severity failure;
	assert RAM(20828) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(20828))))  severity failure;
	assert RAM(20829) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20829))))  severity failure;
	assert RAM(20830) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20830))))  severity failure;
	assert RAM(20831) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20831))))  severity failure;
	assert RAM(20832) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20832))))  severity failure;
	assert RAM(20833) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20833))))  severity failure;
	assert RAM(20834) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20834))))  severity failure;
	assert RAM(20835) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(20835))))  severity failure;
	assert RAM(20836) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20836))))  severity failure;
	assert RAM(20837) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20837))))  severity failure;
	assert RAM(20838) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20838))))  severity failure;
	assert RAM(20839) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20839))))  severity failure;
	assert RAM(20840) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20840))))  severity failure;
	assert RAM(20841) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20841))))  severity failure;
	assert RAM(20842) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20842))))  severity failure;
	assert RAM(20843) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20843))))  severity failure;
	assert RAM(20844) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20844))))  severity failure;
	assert RAM(20845) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20845))))  severity failure;
	assert RAM(20846) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20846))))  severity failure;
	assert RAM(20847) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20847))))  severity failure;
	assert RAM(20848) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20848))))  severity failure;
	assert RAM(20849) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20849))))  severity failure;
	assert RAM(20850) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20850))))  severity failure;
	assert RAM(20851) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20851))))  severity failure;
	assert RAM(20852) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20852))))  severity failure;
	assert RAM(20853) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20853))))  severity failure;
	assert RAM(20854) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20854))))  severity failure;
	assert RAM(20855) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20855))))  severity failure;
	assert RAM(20856) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20856))))  severity failure;
	assert RAM(20857) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(20857))))  severity failure;
	assert RAM(20858) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20858))))  severity failure;
	assert RAM(20859) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20859))))  severity failure;
	assert RAM(20860) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20860))))  severity failure;
	assert RAM(20861) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(20861))))  severity failure;
	assert RAM(20862) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20862))))  severity failure;
	assert RAM(20863) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20863))))  severity failure;
	assert RAM(20864) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20864))))  severity failure;
	assert RAM(20865) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20865))))  severity failure;
	assert RAM(20866) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20866))))  severity failure;
	assert RAM(20867) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20867))))  severity failure;
	assert RAM(20868) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20868))))  severity failure;
	assert RAM(20869) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20869))))  severity failure;
	assert RAM(20870) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(20870))))  severity failure;
	assert RAM(20871) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(20871))))  severity failure;
	assert RAM(20872) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20872))))  severity failure;
	assert RAM(20873) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20873))))  severity failure;
	assert RAM(20874) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20874))))  severity failure;
	assert RAM(20875) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(20875))))  severity failure;
	assert RAM(20876) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20876))))  severity failure;
	assert RAM(20877) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20877))))  severity failure;
	assert RAM(20878) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20878))))  severity failure;
	assert RAM(20879) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20879))))  severity failure;
	assert RAM(20880) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20880))))  severity failure;
	assert RAM(20881) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20881))))  severity failure;
	assert RAM(20882) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20882))))  severity failure;
	assert RAM(20883) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20883))))  severity failure;
	assert RAM(20884) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20884))))  severity failure;
	assert RAM(20885) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20885))))  severity failure;
	assert RAM(20886) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20886))))  severity failure;
	assert RAM(20887) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20887))))  severity failure;
	assert RAM(20888) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20888))))  severity failure;
	assert RAM(20889) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20889))))  severity failure;
	assert RAM(20890) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20890))))  severity failure;
	assert RAM(20891) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20891))))  severity failure;
	assert RAM(20892) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20892))))  severity failure;
	assert RAM(20893) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20893))))  severity failure;
	assert RAM(20894) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20894))))  severity failure;
	assert RAM(20895) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20895))))  severity failure;
	assert RAM(20896) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20896))))  severity failure;
	assert RAM(20897) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20897))))  severity failure;
	assert RAM(20898) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20898))))  severity failure;
	assert RAM(20899) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20899))))  severity failure;
	assert RAM(20900) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20900))))  severity failure;
	assert RAM(20901) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20901))))  severity failure;
	assert RAM(20902) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20902))))  severity failure;
	assert RAM(20903) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20903))))  severity failure;
	assert RAM(20904) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20904))))  severity failure;
	assert RAM(20905) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20905))))  severity failure;
	assert RAM(20906) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20906))))  severity failure;
	assert RAM(20907) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(20907))))  severity failure;
	assert RAM(20908) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20908))))  severity failure;
	assert RAM(20909) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20909))))  severity failure;
	assert RAM(20910) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20910))))  severity failure;
	assert RAM(20911) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20911))))  severity failure;
	assert RAM(20912) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20912))))  severity failure;
	assert RAM(20913) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20913))))  severity failure;
	assert RAM(20914) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20914))))  severity failure;
	assert RAM(20915) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20915))))  severity failure;
	assert RAM(20916) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20916))))  severity failure;
	assert RAM(20917) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20917))))  severity failure;
	assert RAM(20918) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20918))))  severity failure;
	assert RAM(20919) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20919))))  severity failure;
	assert RAM(20920) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20920))))  severity failure;
	assert RAM(20921) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20921))))  severity failure;
	assert RAM(20922) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20922))))  severity failure;
	assert RAM(20923) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20923))))  severity failure;
	assert RAM(20924) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20924))))  severity failure;
	assert RAM(20925) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20925))))  severity failure;
	assert RAM(20926) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(20926))))  severity failure;
	assert RAM(20927) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20927))))  severity failure;
	assert RAM(20928) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20928))))  severity failure;
	assert RAM(20929) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(20929))))  severity failure;
	assert RAM(20930) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20930))))  severity failure;
	assert RAM(20931) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20931))))  severity failure;
	assert RAM(20932) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20932))))  severity failure;
	assert RAM(20933) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20933))))  severity failure;
	assert RAM(20934) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20934))))  severity failure;
	assert RAM(20935) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20935))))  severity failure;
	assert RAM(20936) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20936))))  severity failure;
	assert RAM(20937) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20937))))  severity failure;
	assert RAM(20938) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20938))))  severity failure;
	assert RAM(20939) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(20939))))  severity failure;
	assert RAM(20940) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20940))))  severity failure;
	assert RAM(20941) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20941))))  severity failure;
	assert RAM(20942) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20942))))  severity failure;
	assert RAM(20943) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20943))))  severity failure;
	assert RAM(20944) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20944))))  severity failure;
	assert RAM(20945) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20945))))  severity failure;
	assert RAM(20946) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20946))))  severity failure;
	assert RAM(20947) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20947))))  severity failure;
	assert RAM(20948) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20948))))  severity failure;
	assert RAM(20949) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20949))))  severity failure;
	assert RAM(20950) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20950))))  severity failure;
	assert RAM(20951) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20951))))  severity failure;
	assert RAM(20952) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20952))))  severity failure;
	assert RAM(20953) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20953))))  severity failure;
	assert RAM(20954) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20954))))  severity failure;
	assert RAM(20955) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20955))))  severity failure;
	assert RAM(20956) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20956))))  severity failure;
	assert RAM(20957) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20957))))  severity failure;
	assert RAM(20958) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20958))))  severity failure;
	assert RAM(20959) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20959))))  severity failure;
	assert RAM(20960) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(20960))))  severity failure;
	assert RAM(20961) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(20961))))  severity failure;
	assert RAM(20962) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20962))))  severity failure;
	assert RAM(20963) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20963))))  severity failure;
	assert RAM(20964) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20964))))  severity failure;
	assert RAM(20965) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20965))))  severity failure;
	assert RAM(20966) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20966))))  severity failure;
	assert RAM(20967) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20967))))  severity failure;
	assert RAM(20968) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20968))))  severity failure;
	assert RAM(20969) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20969))))  severity failure;
	assert RAM(20970) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20970))))  severity failure;
	assert RAM(20971) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20971))))  severity failure;
	assert RAM(20972) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20972))))  severity failure;
	assert RAM(20973) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20973))))  severity failure;
	assert RAM(20974) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20974))))  severity failure;
	assert RAM(20975) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20975))))  severity failure;
	assert RAM(20976) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20976))))  severity failure;
	assert RAM(20977) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20977))))  severity failure;
	assert RAM(20978) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20978))))  severity failure;
	assert RAM(20979) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20979))))  severity failure;
	assert RAM(20980) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20980))))  severity failure;
	assert RAM(20981) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20981))))  severity failure;
	assert RAM(20982) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20982))))  severity failure;
	assert RAM(20983) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20983))))  severity failure;
	assert RAM(20984) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(20984))))  severity failure;
	assert RAM(20985) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20985))))  severity failure;
	assert RAM(20986) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20986))))  severity failure;
	assert RAM(20987) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20987))))  severity failure;
	assert RAM(20988) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20988))))  severity failure;
	assert RAM(20989) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20989))))  severity failure;
	assert RAM(20990) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(20990))))  severity failure;
	assert RAM(20991) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20991))))  severity failure;
	assert RAM(20992) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20992))))  severity failure;
	assert RAM(20993) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20993))))  severity failure;
	assert RAM(20994) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20994))))  severity failure;
	assert RAM(20995) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20995))))  severity failure;
	assert RAM(20996) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20996))))  severity failure;
	assert RAM(20997) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20997))))  severity failure;
	assert RAM(20998) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20998))))  severity failure;
	assert RAM(20999) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20999))))  severity failure;
	assert RAM(21000) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(21000))))  severity failure;
	assert RAM(21001) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21001))))  severity failure;
	assert RAM(21002) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21002))))  severity failure;
	assert RAM(21003) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21003))))  severity failure;
	assert RAM(21004) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21004))))  severity failure;
	assert RAM(21005) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21005))))  severity failure;
	assert RAM(21006) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21006))))  severity failure;
	assert RAM(21007) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21007))))  severity failure;
	assert RAM(21008) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21008))))  severity failure;
	assert RAM(21009) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21009))))  severity failure;
	assert RAM(21010) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21010))))  severity failure;
	assert RAM(21011) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21011))))  severity failure;
	assert RAM(21012) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21012))))  severity failure;
	assert RAM(21013) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21013))))  severity failure;
	assert RAM(21014) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21014))))  severity failure;
	assert RAM(21015) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21015))))  severity failure;
	assert RAM(21016) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21016))))  severity failure;
	assert RAM(21017) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21017))))  severity failure;
	assert RAM(21018) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21018))))  severity failure;
	assert RAM(21019) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21019))))  severity failure;
	assert RAM(21020) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21020))))  severity failure;
	assert RAM(21021) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21021))))  severity failure;
	assert RAM(21022) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21022))))  severity failure;
	assert RAM(21023) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(21023))))  severity failure;
	assert RAM(21024) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21024))))  severity failure;
	assert RAM(21025) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21025))))  severity failure;
	assert RAM(21026) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21026))))  severity failure;
	assert RAM(21027) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21027))))  severity failure;
	assert RAM(21028) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21028))))  severity failure;
	assert RAM(21029) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21029))))  severity failure;
	assert RAM(21030) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21030))))  severity failure;
	assert RAM(21031) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21031))))  severity failure;
	assert RAM(21032) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21032))))  severity failure;
	assert RAM(21033) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21033))))  severity failure;
	assert RAM(21034) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21034))))  severity failure;
	assert RAM(21035) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21035))))  severity failure;
	assert RAM(21036) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21036))))  severity failure;
	assert RAM(21037) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21037))))  severity failure;
	assert RAM(21038) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21038))))  severity failure;
	assert RAM(21039) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21039))))  severity failure;
	assert RAM(21040) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21040))))  severity failure;
	assert RAM(21041) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21041))))  severity failure;
	assert RAM(21042) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21042))))  severity failure;
	assert RAM(21043) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21043))))  severity failure;
	assert RAM(21044) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21044))))  severity failure;
	assert RAM(21045) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21045))))  severity failure;
	assert RAM(21046) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21046))))  severity failure;
	assert RAM(21047) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21047))))  severity failure;
	assert RAM(21048) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(21048))))  severity failure;
	assert RAM(21049) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21049))))  severity failure;
	assert RAM(21050) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21050))))  severity failure;
	assert RAM(21051) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21051))))  severity failure;
	assert RAM(21052) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21052))))  severity failure;
	assert RAM(21053) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(21053))))  severity failure;
	assert RAM(21054) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21054))))  severity failure;
	assert RAM(21055) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21055))))  severity failure;
	assert RAM(21056) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(21056))))  severity failure;
	assert RAM(21057) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21057))))  severity failure;
	assert RAM(21058) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21058))))  severity failure;
	assert RAM(21059) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21059))))  severity failure;
	assert RAM(21060) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21060))))  severity failure;
	assert RAM(21061) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21061))))  severity failure;
	assert RAM(21062) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21062))))  severity failure;
	assert RAM(21063) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21063))))  severity failure;
	assert RAM(21064) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(21064))))  severity failure;
	assert RAM(21065) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21065))))  severity failure;
	assert RAM(21066) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21066))))  severity failure;
	assert RAM(21067) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21067))))  severity failure;
	assert RAM(21068) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21068))))  severity failure;
	assert RAM(21069) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21069))))  severity failure;
	assert RAM(21070) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21070))))  severity failure;
	assert RAM(21071) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(21071))))  severity failure;
	assert RAM(21072) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21072))))  severity failure;
	assert RAM(21073) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(21073))))  severity failure;
	assert RAM(21074) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21074))))  severity failure;
	assert RAM(21075) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21075))))  severity failure;
	assert RAM(21076) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21076))))  severity failure;
	assert RAM(21077) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21077))))  severity failure;
	assert RAM(21078) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21078))))  severity failure;
	assert RAM(21079) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(21079))))  severity failure;
	assert RAM(21080) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21080))))  severity failure;
	assert RAM(21081) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21081))))  severity failure;
	assert RAM(21082) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(21082))))  severity failure;
	assert RAM(21083) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21083))))  severity failure;
	assert RAM(21084) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21084))))  severity failure;
	assert RAM(21085) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21085))))  severity failure;
	assert RAM(21086) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21086))))  severity failure;
	assert RAM(21087) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21087))))  severity failure;
	assert RAM(21088) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21088))))  severity failure;
	assert RAM(21089) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21089))))  severity failure;
	assert RAM(21090) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21090))))  severity failure;
	assert RAM(21091) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(21091))))  severity failure;
	assert RAM(21092) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21092))))  severity failure;
	assert RAM(21093) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21093))))  severity failure;
	assert RAM(21094) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21094))))  severity failure;
	assert RAM(21095) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21095))))  severity failure;
	assert RAM(21096) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21096))))  severity failure;
	assert RAM(21097) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21097))))  severity failure;
	assert RAM(21098) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21098))))  severity failure;
	assert RAM(21099) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21099))))  severity failure;
	assert RAM(21100) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21100))))  severity failure;
	assert RAM(21101) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21101))))  severity failure;
	assert RAM(21102) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21102))))  severity failure;
	assert RAM(21103) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21103))))  severity failure;
	assert RAM(21104) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21104))))  severity failure;
	assert RAM(21105) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21105))))  severity failure;
	assert RAM(21106) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21106))))  severity failure;
	assert RAM(21107) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21107))))  severity failure;
	assert RAM(21108) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21108))))  severity failure;
	assert RAM(21109) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21109))))  severity failure;
	assert RAM(21110) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21110))))  severity failure;
	assert RAM(21111) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(21111))))  severity failure;
	assert RAM(21112) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21112))))  severity failure;
	assert RAM(21113) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21113))))  severity failure;
	assert RAM(21114) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21114))))  severity failure;
	assert RAM(21115) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21115))))  severity failure;
	assert RAM(21116) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21116))))  severity failure;
	assert RAM(21117) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21117))))  severity failure;
	assert RAM(21118) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21118))))  severity failure;
	assert RAM(21119) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21119))))  severity failure;
	assert RAM(21120) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21120))))  severity failure;
	assert RAM(21121) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21121))))  severity failure;
	assert RAM(21122) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21122))))  severity failure;
	assert RAM(21123) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21123))))  severity failure;
	assert RAM(21124) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21124))))  severity failure;
	assert RAM(21125) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21125))))  severity failure;
	assert RAM(21126) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21126))))  severity failure;
	assert RAM(21127) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21127))))  severity failure;
	assert RAM(21128) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21128))))  severity failure;
	assert RAM(21129) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21129))))  severity failure;
	assert RAM(21130) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21130))))  severity failure;
	assert RAM(21131) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21131))))  severity failure;
	assert RAM(21132) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21132))))  severity failure;
	assert RAM(21133) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21133))))  severity failure;
	assert RAM(21134) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21134))))  severity failure;
	assert RAM(21135) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21135))))  severity failure;
	assert RAM(21136) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21136))))  severity failure;
	assert RAM(21137) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21137))))  severity failure;
	assert RAM(21138) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21138))))  severity failure;
	assert RAM(21139) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21139))))  severity failure;
	assert RAM(21140) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21140))))  severity failure;
	assert RAM(21141) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21141))))  severity failure;
	assert RAM(21142) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21142))))  severity failure;
	assert RAM(21143) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21143))))  severity failure;
	assert RAM(21144) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21144))))  severity failure;
	assert RAM(21145) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(21145))))  severity failure;
	assert RAM(21146) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21146))))  severity failure;
	assert RAM(21147) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21147))))  severity failure;
	assert RAM(21148) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21148))))  severity failure;
	assert RAM(21149) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21149))))  severity failure;
	assert RAM(21150) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(21150))))  severity failure;
	assert RAM(21151) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21151))))  severity failure;
	assert RAM(21152) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21152))))  severity failure;
	assert RAM(21153) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21153))))  severity failure;
	assert RAM(21154) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21154))))  severity failure;
	assert RAM(21155) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21155))))  severity failure;
	assert RAM(21156) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(21156))))  severity failure;
	assert RAM(21157) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21157))))  severity failure;
	assert RAM(21158) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21158))))  severity failure;
	assert RAM(21159) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21159))))  severity failure;
	assert RAM(21160) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(21160))))  severity failure;
	assert RAM(21161) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21161))))  severity failure;
	assert RAM(21162) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21162))))  severity failure;
	assert RAM(21163) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21163))))  severity failure;
	assert RAM(21164) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21164))))  severity failure;
	assert RAM(21165) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21165))))  severity failure;
	assert RAM(21166) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21166))))  severity failure;
	assert RAM(21167) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21167))))  severity failure;
	assert RAM(21168) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21168))))  severity failure;
	assert RAM(21169) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21169))))  severity failure;
	assert RAM(21170) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21170))))  severity failure;
	assert RAM(21171) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21171))))  severity failure;
	assert RAM(21172) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21172))))  severity failure;
	assert RAM(21173) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21173))))  severity failure;
	assert RAM(21174) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21174))))  severity failure;
	assert RAM(21175) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21175))))  severity failure;
	assert RAM(21176) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21176))))  severity failure;
	assert RAM(21177) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21177))))  severity failure;
	assert RAM(21178) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21178))))  severity failure;
	assert RAM(21179) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(21179))))  severity failure;
	assert RAM(21180) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21180))))  severity failure;
	assert RAM(21181) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21181))))  severity failure;
	assert RAM(21182) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21182))))  severity failure;
	assert RAM(21183) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21183))))  severity failure;
	assert RAM(21184) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21184))))  severity failure;
	assert RAM(21185) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21185))))  severity failure;
	assert RAM(21186) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21186))))  severity failure;
	assert RAM(21187) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21187))))  severity failure;
	assert RAM(21188) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21188))))  severity failure;
	assert RAM(21189) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21189))))  severity failure;
	assert RAM(21190) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21190))))  severity failure;
	assert RAM(21191) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21191))))  severity failure;
	assert RAM(21192) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(21192))))  severity failure;
	assert RAM(21193) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21193))))  severity failure;
	assert RAM(21194) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21194))))  severity failure;
	assert RAM(21195) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21195))))  severity failure;
	assert RAM(21196) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21196))))  severity failure;
	assert RAM(21197) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21197))))  severity failure;
	assert RAM(21198) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21198))))  severity failure;
	assert RAM(21199) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21199))))  severity failure;
	assert RAM(21200) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(21200))))  severity failure;
	assert RAM(21201) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21201))))  severity failure;
	assert RAM(21202) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21202))))  severity failure;
	assert RAM(21203) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(21203))))  severity failure;
	assert RAM(21204) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(21204))))  severity failure;
	assert RAM(21205) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21205))))  severity failure;
	assert RAM(21206) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21206))))  severity failure;
	assert RAM(21207) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21207))))  severity failure;
	assert RAM(21208) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21208))))  severity failure;
	assert RAM(21209) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21209))))  severity failure;
	assert RAM(21210) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21210))))  severity failure;
	assert RAM(21211) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(21211))))  severity failure;
	assert RAM(21212) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(21212))))  severity failure;
	assert RAM(21213) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21213))))  severity failure;
	assert RAM(21214) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21214))))  severity failure;
	assert RAM(21215) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21215))))  severity failure;
	assert RAM(21216) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21216))))  severity failure;
	assert RAM(21217) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21217))))  severity failure;
	assert RAM(21218) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21218))))  severity failure;
	assert RAM(21219) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21219))))  severity failure;
	assert RAM(21220) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21220))))  severity failure;
	assert RAM(21221) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21221))))  severity failure;
	assert RAM(21222) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21222))))  severity failure;
	assert RAM(21223) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21223))))  severity failure;
	assert RAM(21224) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21224))))  severity failure;
	assert RAM(21225) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21225))))  severity failure;
	assert RAM(21226) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21226))))  severity failure;
	assert RAM(21227) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21227))))  severity failure;
	assert RAM(21228) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(21228))))  severity failure;
	assert RAM(21229) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21229))))  severity failure;
	assert RAM(21230) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21230))))  severity failure;
	assert RAM(21231) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21231))))  severity failure;
	assert RAM(21232) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21232))))  severity failure;
	assert RAM(21233) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21233))))  severity failure;
	assert RAM(21234) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21234))))  severity failure;
	assert RAM(21235) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21235))))  severity failure;
	assert RAM(21236) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21236))))  severity failure;
	assert RAM(21237) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21237))))  severity failure;
	assert RAM(21238) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21238))))  severity failure;
	assert RAM(21239) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21239))))  severity failure;
	assert RAM(21240) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21240))))  severity failure;
	assert RAM(21241) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21241))))  severity failure;
	assert RAM(21242) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21242))))  severity failure;
	assert RAM(21243) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21243))))  severity failure;
	assert RAM(21244) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21244))))  severity failure;
	assert RAM(21245) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21245))))  severity failure;
	assert RAM(21246) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21246))))  severity failure;
	assert RAM(21247) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(21247))))  severity failure;
	assert RAM(21248) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21248))))  severity failure;
	assert RAM(21249) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21249))))  severity failure;
	assert RAM(21250) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21250))))  severity failure;
	assert RAM(21251) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21251))))  severity failure;
	assert RAM(21252) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21252))))  severity failure;
	assert RAM(21253) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21253))))  severity failure;
	assert RAM(21254) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21254))))  severity failure;
	assert RAM(21255) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21255))))  severity failure;
	assert RAM(21256) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21256))))  severity failure;
	assert RAM(21257) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(21257))))  severity failure;
	assert RAM(21258) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21258))))  severity failure;
	assert RAM(21259) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21259))))  severity failure;
	assert RAM(21260) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21260))))  severity failure;
	assert RAM(21261) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21261))))  severity failure;
	assert RAM(21262) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21262))))  severity failure;
	assert RAM(21263) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21263))))  severity failure;
	assert RAM(21264) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21264))))  severity failure;
	assert RAM(21265) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21265))))  severity failure;
	assert RAM(21266) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21266))))  severity failure;
	assert RAM(21267) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21267))))  severity failure;
	assert RAM(21268) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21268))))  severity failure;
	assert RAM(21269) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(21269))))  severity failure;
	assert RAM(21270) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(21270))))  severity failure;
	assert RAM(21271) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21271))))  severity failure;
	assert RAM(21272) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21272))))  severity failure;
	assert RAM(21273) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21273))))  severity failure;
	assert RAM(21274) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21274))))  severity failure;
	assert RAM(21275) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21275))))  severity failure;
	assert RAM(21276) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21276))))  severity failure;
	assert RAM(21277) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21277))))  severity failure;
	assert RAM(21278) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21278))))  severity failure;
	assert RAM(21279) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21279))))  severity failure;
	assert RAM(21280) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21280))))  severity failure;
	assert RAM(21281) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21281))))  severity failure;
	assert RAM(21282) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21282))))  severity failure;
	assert RAM(21283) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21283))))  severity failure;
	assert RAM(21284) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21284))))  severity failure;
	assert RAM(21285) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21285))))  severity failure;
	assert RAM(21286) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21286))))  severity failure;
	assert RAM(21287) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21287))))  severity failure;
	assert RAM(21288) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21288))))  severity failure;
	assert RAM(21289) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21289))))  severity failure;
	assert RAM(21290) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(21290))))  severity failure;
	assert RAM(21291) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21291))))  severity failure;
	assert RAM(21292) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(21292))))  severity failure;
	assert RAM(21293) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21293))))  severity failure;
	assert RAM(21294) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21294))))  severity failure;
	assert RAM(21295) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(21295))))  severity failure;
	assert RAM(21296) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21296))))  severity failure;
	assert RAM(21297) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(21297))))  severity failure;
	assert RAM(21298) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21298))))  severity failure;
	assert RAM(21299) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21299))))  severity failure;
	assert RAM(21300) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21300))))  severity failure;
	assert RAM(21301) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21301))))  severity failure;
	assert RAM(21302) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21302))))  severity failure;
	assert RAM(21303) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(21303))))  severity failure;
	assert RAM(21304) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21304))))  severity failure;
	assert RAM(21305) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21305))))  severity failure;
	assert RAM(21306) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21306))))  severity failure;
	assert RAM(21307) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(21307))))  severity failure;
	assert RAM(21308) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21308))))  severity failure;
	assert RAM(21309) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(21309))))  severity failure;
	assert RAM(21310) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21310))))  severity failure;
	assert RAM(21311) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21311))))  severity failure;
	assert RAM(21312) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21312))))  severity failure;
	assert RAM(21313) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21313))))  severity failure;
	assert RAM(21314) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21314))))  severity failure;
	assert RAM(21315) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21315))))  severity failure;
	assert RAM(21316) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21316))))  severity failure;
	assert RAM(21317) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21317))))  severity failure;
	assert RAM(21318) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21318))))  severity failure;
	assert RAM(21319) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21319))))  severity failure;
	assert RAM(21320) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21320))))  severity failure;
	assert RAM(21321) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21321))))  severity failure;
	assert RAM(21322) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21322))))  severity failure;
	assert RAM(21323) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21323))))  severity failure;
	assert RAM(21324) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21324))))  severity failure;
	assert RAM(21325) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21325))))  severity failure;
	assert RAM(21326) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(21326))))  severity failure;
	assert RAM(21327) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21327))))  severity failure;
	assert RAM(21328) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21328))))  severity failure;
	assert RAM(21329) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21329))))  severity failure;
	assert RAM(21330) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21330))))  severity failure;
	assert RAM(21331) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21331))))  severity failure;
	assert RAM(21332) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(21332))))  severity failure;
	assert RAM(21333) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21333))))  severity failure;
	assert RAM(21334) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21334))))  severity failure;
	assert RAM(21335) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21335))))  severity failure;
	assert RAM(21336) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21336))))  severity failure;
	assert RAM(21337) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21337))))  severity failure;
	assert RAM(21338) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21338))))  severity failure;
	assert RAM(21339) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21339))))  severity failure;
	assert RAM(21340) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21340))))  severity failure;
	assert RAM(21341) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21341))))  severity failure;
	assert RAM(21342) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21342))))  severity failure;
	assert RAM(21343) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21343))))  severity failure;
	assert RAM(21344) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21344))))  severity failure;
	assert RAM(21345) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21345))))  severity failure;
	assert RAM(21346) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21346))))  severity failure;
	assert RAM(21347) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(21347))))  severity failure;
	assert RAM(21348) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21348))))  severity failure;
	assert RAM(21349) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21349))))  severity failure;
	assert RAM(21350) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21350))))  severity failure;
	assert RAM(21351) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21351))))  severity failure;
	assert RAM(21352) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21352))))  severity failure;
	assert RAM(21353) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(21353))))  severity failure;
	assert RAM(21354) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21354))))  severity failure;
	assert RAM(21355) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21355))))  severity failure;
	assert RAM(21356) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21356))))  severity failure;
	assert RAM(21357) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21357))))  severity failure;
	assert RAM(21358) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21358))))  severity failure;
	assert RAM(21359) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(21359))))  severity failure;
	assert RAM(21360) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21360))))  severity failure;
	assert RAM(21361) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21361))))  severity failure;
	assert RAM(21362) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21362))))  severity failure;
	assert RAM(21363) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21363))))  severity failure;
	assert RAM(21364) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21364))))  severity failure;
	assert RAM(21365) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21365))))  severity failure;
	assert RAM(21366) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21366))))  severity failure;
	assert RAM(21367) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21367))))  severity failure;
	assert RAM(21368) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21368))))  severity failure;
	assert RAM(21369) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21369))))  severity failure;
	assert RAM(21370) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21370))))  severity failure;
	assert RAM(21371) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(21371))))  severity failure;
	assert RAM(21372) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21372))))  severity failure;
	assert RAM(21373) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21373))))  severity failure;
	assert RAM(21374) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21374))))  severity failure;
	assert RAM(21375) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21375))))  severity failure;
	assert RAM(21376) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21376))))  severity failure;
	assert RAM(21377) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21377))))  severity failure;
	assert RAM(21378) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21378))))  severity failure;
	assert RAM(21379) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21379))))  severity failure;
	assert RAM(21380) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21380))))  severity failure;
	assert RAM(21381) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21381))))  severity failure;
	assert RAM(21382) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21382))))  severity failure;
	assert RAM(21383) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21383))))  severity failure;
	assert RAM(21384) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(21384))))  severity failure;
	assert RAM(21385) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21385))))  severity failure;
	assert RAM(21386) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(21386))))  severity failure;
	assert RAM(21387) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21387))))  severity failure;
	assert RAM(21388) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21388))))  severity failure;
	assert RAM(21389) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21389))))  severity failure;
	assert RAM(21390) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21390))))  severity failure;
	assert RAM(21391) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21391))))  severity failure;
	assert RAM(21392) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21392))))  severity failure;
	assert RAM(21393) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21393))))  severity failure;
	assert RAM(21394) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21394))))  severity failure;
	assert RAM(21395) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21395))))  severity failure;
	assert RAM(21396) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21396))))  severity failure;
	assert RAM(21397) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21397))))  severity failure;
	assert RAM(21398) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21398))))  severity failure;
	assert RAM(21399) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(21399))))  severity failure;
	assert RAM(21400) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21400))))  severity failure;
	assert RAM(21401) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21401))))  severity failure;
	assert RAM(21402) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(21402))))  severity failure;
	assert RAM(21403) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21403))))  severity failure;
	assert RAM(21404) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(21404))))  severity failure;
	assert RAM(21405) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21405))))  severity failure;
	assert RAM(21406) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21406))))  severity failure;
	assert RAM(21407) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21407))))  severity failure;
	assert RAM(21408) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21408))))  severity failure;
	assert RAM(21409) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21409))))  severity failure;
	assert RAM(21410) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21410))))  severity failure;
	assert RAM(21411) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21411))))  severity failure;
	assert RAM(21412) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21412))))  severity failure;
	assert RAM(21413) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21413))))  severity failure;
	assert RAM(21414) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21414))))  severity failure;
	assert RAM(21415) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21415))))  severity failure;
	assert RAM(21416) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21416))))  severity failure;
	assert RAM(21417) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21417))))  severity failure;
	assert RAM(21418) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21418))))  severity failure;
	assert RAM(21419) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21419))))  severity failure;
	assert RAM(21420) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21420))))  severity failure;
	assert RAM(21421) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21421))))  severity failure;
	assert RAM(21422) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21422))))  severity failure;
	assert RAM(21423) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21423))))  severity failure;
	assert RAM(21424) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21424))))  severity failure;
	assert RAM(21425) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21425))))  severity failure;
	assert RAM(21426) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21426))))  severity failure;
	assert RAM(21427) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21427))))  severity failure;
	assert RAM(21428) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21428))))  severity failure;
	assert RAM(21429) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(21429))))  severity failure;
	assert RAM(21430) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21430))))  severity failure;
	assert RAM(21431) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21431))))  severity failure;
	assert RAM(21432) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(21432))))  severity failure;
	assert RAM(21433) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21433))))  severity failure;
	assert RAM(21434) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21434))))  severity failure;
	assert RAM(21435) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21435))))  severity failure;
	assert RAM(21436) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21436))))  severity failure;
	assert RAM(21437) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21437))))  severity failure;
	assert RAM(21438) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(21438))))  severity failure;
	assert RAM(21439) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21439))))  severity failure;
	assert RAM(21440) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21440))))  severity failure;
	assert RAM(21441) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(21441))))  severity failure;
	assert RAM(21442) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(21442))))  severity failure;
	assert RAM(21443) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21443))))  severity failure;
	assert RAM(21444) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21444))))  severity failure;
	assert RAM(21445) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21445))))  severity failure;
	assert RAM(21446) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(21446))))  severity failure;
	assert RAM(21447) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(21447))))  severity failure;
	assert RAM(21448) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21448))))  severity failure;
	assert RAM(21449) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21449))))  severity failure;
	assert RAM(21450) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21450))))  severity failure;
	assert RAM(21451) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(21451))))  severity failure;
	assert RAM(21452) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21452))))  severity failure;
	assert RAM(21453) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21453))))  severity failure;
	assert RAM(21454) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21454))))  severity failure;
	assert RAM(21455) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21455))))  severity failure;
	assert RAM(21456) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21456))))  severity failure;
	assert RAM(21457) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21457))))  severity failure;
	assert RAM(21458) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21458))))  severity failure;
	assert RAM(21459) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21459))))  severity failure;
	assert RAM(21460) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(21460))))  severity failure;
	assert RAM(21461) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21461))))  severity failure;
	assert RAM(21462) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21462))))  severity failure;
	assert RAM(21463) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21463))))  severity failure;
	assert RAM(21464) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21464))))  severity failure;
	assert RAM(21465) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21465))))  severity failure;
	assert RAM(21466) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21466))))  severity failure;
	assert RAM(21467) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21467))))  severity failure;
	assert RAM(21468) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21468))))  severity failure;
	assert RAM(21469) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21469))))  severity failure;
	assert RAM(21470) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(21470))))  severity failure;
	assert RAM(21471) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(21471))))  severity failure;
	assert RAM(21472) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21472))))  severity failure;
	assert RAM(21473) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21473))))  severity failure;
	assert RAM(21474) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21474))))  severity failure;
	assert RAM(21475) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21475))))  severity failure;
	assert RAM(21476) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21476))))  severity failure;
	assert RAM(21477) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21477))))  severity failure;
	assert RAM(21478) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21478))))  severity failure;
	assert RAM(21479) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21479))))  severity failure;
	assert RAM(21480) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21480))))  severity failure;
	assert RAM(21481) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21481))))  severity failure;
	assert RAM(21482) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21482))))  severity failure;
	assert RAM(21483) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21483))))  severity failure;
	assert RAM(21484) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(21484))))  severity failure;
	assert RAM(21485) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21485))))  severity failure;
	assert RAM(21486) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21486))))  severity failure;
	assert RAM(21487) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21487))))  severity failure;
	assert RAM(21488) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21488))))  severity failure;
	assert RAM(21489) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21489))))  severity failure;
	assert RAM(21490) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21490))))  severity failure;
	assert RAM(21491) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21491))))  severity failure;
	assert RAM(21492) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(21492))))  severity failure;
	assert RAM(21493) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21493))))  severity failure;
	assert RAM(21494) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21494))))  severity failure;
	assert RAM(21495) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(21495))))  severity failure;
	assert RAM(21496) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21496))))  severity failure;
	assert RAM(21497) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21497))))  severity failure;
	assert RAM(21498) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21498))))  severity failure;
	assert RAM(21499) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21499))))  severity failure;
	assert RAM(21500) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21500))))  severity failure;
	assert RAM(21501) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21501))))  severity failure;
	assert RAM(21502) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21502))))  severity failure;
	assert RAM(21503) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21503))))  severity failure;
	assert RAM(21504) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21504))))  severity failure;
	assert RAM(21505) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21505))))  severity failure;
	assert RAM(21506) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21506))))  severity failure;
	assert RAM(21507) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21507))))  severity failure;
	assert RAM(21508) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21508))))  severity failure;
	assert RAM(21509) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21509))))  severity failure;
	assert RAM(21510) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21510))))  severity failure;
	assert RAM(21511) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21511))))  severity failure;
	assert RAM(21512) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21512))))  severity failure;
	assert RAM(21513) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21513))))  severity failure;
	assert RAM(21514) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21514))))  severity failure;
	assert RAM(21515) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21515))))  severity failure;
	assert RAM(21516) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21516))))  severity failure;
	assert RAM(21517) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21517))))  severity failure;
	assert RAM(21518) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21518))))  severity failure;
	assert RAM(21519) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21519))))  severity failure;
	assert RAM(21520) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21520))))  severity failure;
	assert RAM(21521) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21521))))  severity failure;
	assert RAM(21522) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21522))))  severity failure;
	assert RAM(21523) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21523))))  severity failure;
	assert RAM(21524) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21524))))  severity failure;
	assert RAM(21525) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21525))))  severity failure;
	assert RAM(21526) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21526))))  severity failure;
	assert RAM(21527) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21527))))  severity failure;
	assert RAM(21528) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21528))))  severity failure;
	assert RAM(21529) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21529))))  severity failure;
	assert RAM(21530) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21530))))  severity failure;
	assert RAM(21531) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21531))))  severity failure;
	assert RAM(21532) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21532))))  severity failure;
	assert RAM(21533) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21533))))  severity failure;
	assert RAM(21534) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21534))))  severity failure;
	assert RAM(21535) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21535))))  severity failure;
	assert RAM(21536) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21536))))  severity failure;
	assert RAM(21537) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21537))))  severity failure;
	assert RAM(21538) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21538))))  severity failure;
	assert RAM(21539) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21539))))  severity failure;
	assert RAM(21540) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21540))))  severity failure;
	assert RAM(21541) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21541))))  severity failure;
	assert RAM(21542) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21542))))  severity failure;
	assert RAM(21543) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21543))))  severity failure;
	assert RAM(21544) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21544))))  severity failure;
	assert RAM(21545) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21545))))  severity failure;
	assert RAM(21546) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21546))))  severity failure;
	assert RAM(21547) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(21547))))  severity failure;
	assert RAM(21548) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21548))))  severity failure;
	assert RAM(21549) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(21549))))  severity failure;
	assert RAM(21550) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21550))))  severity failure;
	assert RAM(21551) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(21551))))  severity failure;
	assert RAM(21552) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21552))))  severity failure;
	assert RAM(21553) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21553))))  severity failure;
	assert RAM(21554) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21554))))  severity failure;
	assert RAM(21555) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(21555))))  severity failure;
	assert RAM(21556) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21556))))  severity failure;
	assert RAM(21557) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21557))))  severity failure;
	assert RAM(21558) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21558))))  severity failure;
	assert RAM(21559) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21559))))  severity failure;
	assert RAM(21560) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21560))))  severity failure;
	assert RAM(21561) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21561))))  severity failure;
	assert RAM(21562) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21562))))  severity failure;
	assert RAM(21563) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(21563))))  severity failure;
	assert RAM(21564) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21564))))  severity failure;
	assert RAM(21565) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21565))))  severity failure;
	assert RAM(21566) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21566))))  severity failure;
	assert RAM(21567) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21567))))  severity failure;
	assert RAM(21568) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21568))))  severity failure;
	assert RAM(21569) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21569))))  severity failure;
	assert RAM(21570) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21570))))  severity failure;
	assert RAM(21571) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21571))))  severity failure;
	assert RAM(21572) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21572))))  severity failure;
	assert RAM(21573) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21573))))  severity failure;
	assert RAM(21574) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21574))))  severity failure;
	assert RAM(21575) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21575))))  severity failure;
	assert RAM(21576) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21576))))  severity failure;
	assert RAM(21577) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21577))))  severity failure;
	assert RAM(21578) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21578))))  severity failure;
	assert RAM(21579) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21579))))  severity failure;
	assert RAM(21580) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(21580))))  severity failure;
	assert RAM(21581) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21581))))  severity failure;
	assert RAM(21582) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21582))))  severity failure;
	assert RAM(21583) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21583))))  severity failure;
	assert RAM(21584) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21584))))  severity failure;
	assert RAM(21585) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21585))))  severity failure;
	assert RAM(21586) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21586))))  severity failure;
	assert RAM(21587) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21587))))  severity failure;
	assert RAM(21588) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(21588))))  severity failure;
	assert RAM(21589) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21589))))  severity failure;
	assert RAM(21590) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21590))))  severity failure;
	assert RAM(21591) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21591))))  severity failure;
	assert RAM(21592) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21592))))  severity failure;
	assert RAM(21593) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(21593))))  severity failure;
	assert RAM(21594) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21594))))  severity failure;
	assert RAM(21595) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21595))))  severity failure;
	assert RAM(21596) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21596))))  severity failure;
	assert RAM(21597) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(21597))))  severity failure;
	assert RAM(21598) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21598))))  severity failure;
	assert RAM(21599) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21599))))  severity failure;
	assert RAM(21600) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21600))))  severity failure;
	assert RAM(21601) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21601))))  severity failure;
	assert RAM(21602) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21602))))  severity failure;
	assert RAM(21603) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21603))))  severity failure;
	assert RAM(21604) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21604))))  severity failure;
	assert RAM(21605) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21605))))  severity failure;
	assert RAM(21606) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(21606))))  severity failure;
	assert RAM(21607) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21607))))  severity failure;
	assert RAM(21608) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21608))))  severity failure;
	assert RAM(21609) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21609))))  severity failure;
	assert RAM(21610) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21610))))  severity failure;
	assert RAM(21611) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(21611))))  severity failure;
	assert RAM(21612) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21612))))  severity failure;
	assert RAM(21613) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21613))))  severity failure;
	assert RAM(21614) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21614))))  severity failure;
	assert RAM(21615) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21615))))  severity failure;
	assert RAM(21616) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21616))))  severity failure;
	assert RAM(21617) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21617))))  severity failure;
	assert RAM(21618) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21618))))  severity failure;
	assert RAM(21619) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21619))))  severity failure;
	assert RAM(21620) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21620))))  severity failure;
	assert RAM(21621) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21621))))  severity failure;
	assert RAM(21622) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21622))))  severity failure;
	assert RAM(21623) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21623))))  severity failure;
	assert RAM(21624) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21624))))  severity failure;
	assert RAM(21625) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21625))))  severity failure;
	assert RAM(21626) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21626))))  severity failure;
	assert RAM(21627) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21627))))  severity failure;
	assert RAM(21628) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21628))))  severity failure;
	assert RAM(21629) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21629))))  severity failure;
	assert RAM(21630) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21630))))  severity failure;
	assert RAM(21631) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21631))))  severity failure;
	assert RAM(21632) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21632))))  severity failure;
	assert RAM(21633) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21633))))  severity failure;
	assert RAM(21634) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21634))))  severity failure;
	assert RAM(21635) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21635))))  severity failure;
	assert RAM(21636) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21636))))  severity failure;
	assert RAM(21637) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21637))))  severity failure;
	assert RAM(21638) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21638))))  severity failure;
	assert RAM(21639) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21639))))  severity failure;
	assert RAM(21640) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21640))))  severity failure;
	assert RAM(21641) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21641))))  severity failure;
	assert RAM(21642) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21642))))  severity failure;
	assert RAM(21643) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21643))))  severity failure;
	assert RAM(21644) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(21644))))  severity failure;
	assert RAM(21645) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21645))))  severity failure;
	assert RAM(21646) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21646))))  severity failure;
	assert RAM(21647) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21647))))  severity failure;
	assert RAM(21648) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(21648))))  severity failure;
	assert RAM(21649) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21649))))  severity failure;
	assert RAM(21650) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21650))))  severity failure;
	assert RAM(21651) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21651))))  severity failure;
	assert RAM(21652) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21652))))  severity failure;
	assert RAM(21653) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21653))))  severity failure;
	assert RAM(21654) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21654))))  severity failure;
	assert RAM(21655) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21655))))  severity failure;
	assert RAM(21656) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21656))))  severity failure;
	assert RAM(21657) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21657))))  severity failure;
	assert RAM(21658) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21658))))  severity failure;
	assert RAM(21659) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21659))))  severity failure;
	assert RAM(21660) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21660))))  severity failure;
	assert RAM(21661) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21661))))  severity failure;
	assert RAM(21662) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(21662))))  severity failure;
	assert RAM(21663) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(21663))))  severity failure;
	assert RAM(21664) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21664))))  severity failure;
	assert RAM(21665) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21665))))  severity failure;
	assert RAM(21666) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21666))))  severity failure;
	assert RAM(21667) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21667))))  severity failure;
	assert RAM(21668) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21668))))  severity failure;
	assert RAM(21669) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21669))))  severity failure;
	assert RAM(21670) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21670))))  severity failure;
	assert RAM(21671) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21671))))  severity failure;
	assert RAM(21672) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21672))))  severity failure;
	assert RAM(21673) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21673))))  severity failure;
	assert RAM(21674) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21674))))  severity failure;
	assert RAM(21675) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21675))))  severity failure;
	assert RAM(21676) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(21676))))  severity failure;
	assert RAM(21677) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(21677))))  severity failure;
	assert RAM(21678) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21678))))  severity failure;
	assert RAM(21679) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21679))))  severity failure;
	assert RAM(21680) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21680))))  severity failure;
	assert RAM(21681) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21681))))  severity failure;
	assert RAM(21682) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(21682))))  severity failure;
	assert RAM(21683) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21683))))  severity failure;
	assert RAM(21684) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21684))))  severity failure;
	assert RAM(21685) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21685))))  severity failure;
	assert RAM(21686) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(21686))))  severity failure;
	assert RAM(21687) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21687))))  severity failure;
	assert RAM(21688) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21688))))  severity failure;
	assert RAM(21689) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21689))))  severity failure;
	assert RAM(21690) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21690))))  severity failure;
	assert RAM(21691) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21691))))  severity failure;
	assert RAM(21692) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21692))))  severity failure;
	assert RAM(21693) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(21693))))  severity failure;
	assert RAM(21694) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21694))))  severity failure;
	assert RAM(21695) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21695))))  severity failure;
	assert RAM(21696) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(21696))))  severity failure;
	assert RAM(21697) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21697))))  severity failure;
	assert RAM(21698) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21698))))  severity failure;
	assert RAM(21699) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(21699))))  severity failure;
	assert RAM(21700) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21700))))  severity failure;
	assert RAM(21701) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21701))))  severity failure;
	assert RAM(21702) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21702))))  severity failure;
	assert RAM(21703) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21703))))  severity failure;
	assert RAM(21704) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21704))))  severity failure;
	assert RAM(21705) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21705))))  severity failure;
	assert RAM(21706) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(21706))))  severity failure;
	assert RAM(21707) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(21707))))  severity failure;
	assert RAM(21708) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21708))))  severity failure;
	assert RAM(21709) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21709))))  severity failure;
	assert RAM(21710) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21710))))  severity failure;
	assert RAM(21711) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21711))))  severity failure;
	assert RAM(21712) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(21712))))  severity failure;
	assert RAM(21713) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21713))))  severity failure;
	assert RAM(21714) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21714))))  severity failure;
	assert RAM(21715) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21715))))  severity failure;
	assert RAM(21716) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21716))))  severity failure;
	assert RAM(21717) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(21717))))  severity failure;
	assert RAM(21718) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21718))))  severity failure;
	assert RAM(21719) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21719))))  severity failure;
	assert RAM(21720) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21720))))  severity failure;
	assert RAM(21721) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21721))))  severity failure;
	assert RAM(21722) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21722))))  severity failure;
	assert RAM(21723) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21723))))  severity failure;
	assert RAM(21724) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21724))))  severity failure;
	assert RAM(21725) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21725))))  severity failure;
	assert RAM(21726) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21726))))  severity failure;
	assert RAM(21727) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21727))))  severity failure;
	assert RAM(21728) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21728))))  severity failure;
	assert RAM(21729) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(21729))))  severity failure;
	assert RAM(21730) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21730))))  severity failure;
	assert RAM(21731) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21731))))  severity failure;
	assert RAM(21732) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21732))))  severity failure;
	assert RAM(21733) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21733))))  severity failure;
	assert RAM(21734) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(21734))))  severity failure;
	assert RAM(21735) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21735))))  severity failure;
	assert RAM(21736) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21736))))  severity failure;
	assert RAM(21737) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21737))))  severity failure;
	assert RAM(21738) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21738))))  severity failure;
	assert RAM(21739) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21739))))  severity failure;
	assert RAM(21740) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21740))))  severity failure;
	assert RAM(21741) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21741))))  severity failure;
	assert RAM(21742) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21742))))  severity failure;
	assert RAM(21743) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21743))))  severity failure;
	assert RAM(21744) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21744))))  severity failure;
	assert RAM(21745) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21745))))  severity failure;
	assert RAM(21746) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21746))))  severity failure;
	assert RAM(21747) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21747))))  severity failure;
	assert RAM(21748) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21748))))  severity failure;
	assert RAM(21749) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21749))))  severity failure;
	assert RAM(21750) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21750))))  severity failure;
	assert RAM(21751) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21751))))  severity failure;
	assert RAM(21752) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21752))))  severity failure;
	assert RAM(21753) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21753))))  severity failure;
	assert RAM(21754) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21754))))  severity failure;
	assert RAM(21755) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21755))))  severity failure;
	assert RAM(21756) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21756))))  severity failure;
	assert RAM(21757) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(21757))))  severity failure;
	assert RAM(21758) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21758))))  severity failure;
	assert RAM(21759) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21759))))  severity failure;
	assert RAM(21760) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21760))))  severity failure;
	assert RAM(21761) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21761))))  severity failure;
	assert RAM(21762) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21762))))  severity failure;
	assert RAM(21763) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21763))))  severity failure;
	assert RAM(21764) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21764))))  severity failure;
	assert RAM(21765) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21765))))  severity failure;
	assert RAM(21766) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21766))))  severity failure;
	assert RAM(21767) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21767))))  severity failure;
	assert RAM(21768) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21768))))  severity failure;
	assert RAM(21769) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21769))))  severity failure;
	assert RAM(21770) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21770))))  severity failure;
	assert RAM(21771) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21771))))  severity failure;
	assert RAM(21772) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21772))))  severity failure;
	assert RAM(21773) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21773))))  severity failure;
	assert RAM(21774) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21774))))  severity failure;
	assert RAM(21775) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21775))))  severity failure;
	assert RAM(21776) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21776))))  severity failure;
	assert RAM(21777) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21777))))  severity failure;
	assert RAM(21778) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21778))))  severity failure;
	assert RAM(21779) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21779))))  severity failure;
	assert RAM(21780) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21780))))  severity failure;
	assert RAM(21781) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21781))))  severity failure;
	assert RAM(21782) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21782))))  severity failure;
	assert RAM(21783) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(21783))))  severity failure;
	assert RAM(21784) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21784))))  severity failure;
	assert RAM(21785) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21785))))  severity failure;
	assert RAM(21786) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21786))))  severity failure;
	assert RAM(21787) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21787))))  severity failure;
	assert RAM(21788) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21788))))  severity failure;
	assert RAM(21789) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(21789))))  severity failure;
	assert RAM(21790) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21790))))  severity failure;
	assert RAM(21791) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21791))))  severity failure;
	assert RAM(21792) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(21792))))  severity failure;
	assert RAM(21793) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21793))))  severity failure;
	assert RAM(21794) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21794))))  severity failure;
	assert RAM(21795) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21795))))  severity failure;
	assert RAM(21796) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21796))))  severity failure;
	assert RAM(21797) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21797))))  severity failure;
	assert RAM(21798) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21798))))  severity failure;
	assert RAM(21799) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21799))))  severity failure;
	assert RAM(21800) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21800))))  severity failure;
	assert RAM(21801) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21801))))  severity failure;
	assert RAM(21802) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21802))))  severity failure;
	assert RAM(21803) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(21803))))  severity failure;
	assert RAM(21804) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21804))))  severity failure;
	assert RAM(21805) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(21805))))  severity failure;
	assert RAM(21806) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(21806))))  severity failure;
	assert RAM(21807) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21807))))  severity failure;
	assert RAM(21808) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21808))))  severity failure;
	assert RAM(21809) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21809))))  severity failure;
	assert RAM(21810) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21810))))  severity failure;
	assert RAM(21811) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21811))))  severity failure;
	assert RAM(21812) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21812))))  severity failure;
	assert RAM(21813) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21813))))  severity failure;
	assert RAM(21814) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21814))))  severity failure;
	assert RAM(21815) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21815))))  severity failure;
	assert RAM(21816) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21816))))  severity failure;
	assert RAM(21817) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21817))))  severity failure;
	assert RAM(21818) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21818))))  severity failure;
	assert RAM(21819) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21819))))  severity failure;
	assert RAM(21820) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21820))))  severity failure;
	assert RAM(21821) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21821))))  severity failure;
	assert RAM(21822) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21822))))  severity failure;
	assert RAM(21823) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21823))))  severity failure;
	assert RAM(21824) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(21824))))  severity failure;
	assert RAM(21825) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21825))))  severity failure;
	assert RAM(21826) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21826))))  severity failure;
	assert RAM(21827) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21827))))  severity failure;
	assert RAM(21828) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21828))))  severity failure;
	assert RAM(21829) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21829))))  severity failure;
	assert RAM(21830) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21830))))  severity failure;
	assert RAM(21831) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21831))))  severity failure;
	assert RAM(21832) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21832))))  severity failure;
	assert RAM(21833) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21833))))  severity failure;
	assert RAM(21834) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21834))))  severity failure;
	assert RAM(21835) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21835))))  severity failure;
	assert RAM(21836) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21836))))  severity failure;
	assert RAM(21837) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21837))))  severity failure;
	assert RAM(21838) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21838))))  severity failure;
	assert RAM(21839) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21839))))  severity failure;
	assert RAM(21840) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(21840))))  severity failure;
	assert RAM(21841) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21841))))  severity failure;
	assert RAM(21842) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21842))))  severity failure;
	assert RAM(21843) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21843))))  severity failure;
	assert RAM(21844) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21844))))  severity failure;
	assert RAM(21845) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21845))))  severity failure;
	assert RAM(21846) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21846))))  severity failure;
	assert RAM(21847) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21847))))  severity failure;
	assert RAM(21848) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21848))))  severity failure;
	assert RAM(21849) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21849))))  severity failure;
	assert RAM(21850) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21850))))  severity failure;
	assert RAM(21851) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21851))))  severity failure;
	assert RAM(21852) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(21852))))  severity failure;
	assert RAM(21853) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21853))))  severity failure;
	assert RAM(21854) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21854))))  severity failure;
	assert RAM(21855) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21855))))  severity failure;
	assert RAM(21856) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21856))))  severity failure;
	assert RAM(21857) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21857))))  severity failure;
	assert RAM(21858) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21858))))  severity failure;
	assert RAM(21859) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21859))))  severity failure;
	assert RAM(21860) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21860))))  severity failure;
	assert RAM(21861) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21861))))  severity failure;
	assert RAM(21862) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21862))))  severity failure;
	assert RAM(21863) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21863))))  severity failure;
	assert RAM(21864) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21864))))  severity failure;
	assert RAM(21865) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21865))))  severity failure;
	assert RAM(21866) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21866))))  severity failure;
	assert RAM(21867) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21867))))  severity failure;
	assert RAM(21868) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21868))))  severity failure;
	assert RAM(21869) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21869))))  severity failure;
	assert RAM(21870) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21870))))  severity failure;
	assert RAM(21871) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21871))))  severity failure;
	assert RAM(21872) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21872))))  severity failure;
	assert RAM(21873) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21873))))  severity failure;
	assert RAM(21874) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21874))))  severity failure;
	assert RAM(21875) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21875))))  severity failure;
	assert RAM(21876) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21876))))  severity failure;
	assert RAM(21877) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21877))))  severity failure;
	assert RAM(21878) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21878))))  severity failure;
	assert RAM(21879) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21879))))  severity failure;
	assert RAM(21880) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21880))))  severity failure;
	assert RAM(21881) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21881))))  severity failure;
	assert RAM(21882) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(21882))))  severity failure;
	assert RAM(21883) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21883))))  severity failure;
	assert RAM(21884) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21884))))  severity failure;
	assert RAM(21885) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(21885))))  severity failure;
	assert RAM(21886) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21886))))  severity failure;
	assert RAM(21887) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21887))))  severity failure;
	assert RAM(21888) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21888))))  severity failure;
	assert RAM(21889) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21889))))  severity failure;
	assert RAM(21890) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21890))))  severity failure;
	assert RAM(21891) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21891))))  severity failure;
	assert RAM(21892) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21892))))  severity failure;
	assert RAM(21893) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21893))))  severity failure;
	assert RAM(21894) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21894))))  severity failure;
	assert RAM(21895) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21895))))  severity failure;
	assert RAM(21896) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21896))))  severity failure;
	assert RAM(21897) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21897))))  severity failure;
	assert RAM(21898) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21898))))  severity failure;
	assert RAM(21899) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21899))))  severity failure;
	assert RAM(21900) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21900))))  severity failure;
	assert RAM(21901) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21901))))  severity failure;
	assert RAM(21902) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21902))))  severity failure;
	assert RAM(21903) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21903))))  severity failure;
	assert RAM(21904) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21904))))  severity failure;
	assert RAM(21905) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21905))))  severity failure;
	assert RAM(21906) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21906))))  severity failure;
	assert RAM(21907) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21907))))  severity failure;
	assert RAM(21908) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21908))))  severity failure;
	assert RAM(21909) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21909))))  severity failure;
	assert RAM(21910) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21910))))  severity failure;
	assert RAM(21911) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(21911))))  severity failure;
	assert RAM(21912) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21912))))  severity failure;
	assert RAM(21913) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21913))))  severity failure;
	assert RAM(21914) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21914))))  severity failure;
	assert RAM(21915) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21915))))  severity failure;
	assert RAM(21916) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21916))))  severity failure;
	assert RAM(21917) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21917))))  severity failure;
	assert RAM(21918) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21918))))  severity failure;
	assert RAM(21919) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(21919))))  severity failure;
	assert RAM(21920) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21920))))  severity failure;
	assert RAM(21921) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21921))))  severity failure;
	assert RAM(21922) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21922))))  severity failure;
	assert RAM(21923) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21923))))  severity failure;
	assert RAM(21924) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21924))))  severity failure;
	assert RAM(21925) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21925))))  severity failure;
	assert RAM(21926) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21926))))  severity failure;
	assert RAM(21927) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21927))))  severity failure;
	assert RAM(21928) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21928))))  severity failure;
	assert RAM(21929) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21929))))  severity failure;
	assert RAM(21930) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21930))))  severity failure;
	assert RAM(21931) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(21931))))  severity failure;
	assert RAM(21932) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21932))))  severity failure;
	assert RAM(21933) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21933))))  severity failure;
	assert RAM(21934) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21934))))  severity failure;
	assert RAM(21935) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21935))))  severity failure;
	assert RAM(21936) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21936))))  severity failure;
	assert RAM(21937) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21937))))  severity failure;
	assert RAM(21938) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21938))))  severity failure;
	assert RAM(21939) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21939))))  severity failure;
	assert RAM(21940) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21940))))  severity failure;
	assert RAM(21941) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21941))))  severity failure;
	assert RAM(21942) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21942))))  severity failure;
	assert RAM(21943) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21943))))  severity failure;
	assert RAM(21944) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21944))))  severity failure;
	assert RAM(21945) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21945))))  severity failure;
	assert RAM(21946) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21946))))  severity failure;
	assert RAM(21947) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(21947))))  severity failure;
	assert RAM(21948) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21948))))  severity failure;
	assert RAM(21949) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21949))))  severity failure;
	assert RAM(21950) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21950))))  severity failure;
	assert RAM(21951) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21951))))  severity failure;
	assert RAM(21952) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21952))))  severity failure;
	assert RAM(21953) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21953))))  severity failure;
	assert RAM(21954) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21954))))  severity failure;
	assert RAM(21955) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21955))))  severity failure;
	assert RAM(21956) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21956))))  severity failure;
	assert RAM(21957) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21957))))  severity failure;
	assert RAM(21958) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21958))))  severity failure;
	assert RAM(21959) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21959))))  severity failure;
	assert RAM(21960) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21960))))  severity failure;
	assert RAM(21961) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21961))))  severity failure;
	assert RAM(21962) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21962))))  severity failure;
	assert RAM(21963) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(21963))))  severity failure;
	assert RAM(21964) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21964))))  severity failure;
	assert RAM(21965) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21965))))  severity failure;
	assert RAM(21966) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21966))))  severity failure;
	assert RAM(21967) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21967))))  severity failure;
	assert RAM(21968) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21968))))  severity failure;
	assert RAM(21969) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21969))))  severity failure;
	assert RAM(21970) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21970))))  severity failure;
	assert RAM(21971) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21971))))  severity failure;
	assert RAM(21972) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21972))))  severity failure;
	assert RAM(21973) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21973))))  severity failure;
	assert RAM(21974) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21974))))  severity failure;
	assert RAM(21975) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21975))))  severity failure;
	assert RAM(21976) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21976))))  severity failure;
	assert RAM(21977) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21977))))  severity failure;
	assert RAM(21978) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21978))))  severity failure;
	assert RAM(21979) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(21979))))  severity failure;
	assert RAM(21980) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21980))))  severity failure;
	assert RAM(21981) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21981))))  severity failure;
	assert RAM(21982) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21982))))  severity failure;
	assert RAM(21983) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21983))))  severity failure;
	assert RAM(21984) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21984))))  severity failure;
	assert RAM(21985) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21985))))  severity failure;
	assert RAM(21986) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21986))))  severity failure;
	assert RAM(21987) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21987))))  severity failure;
	assert RAM(21988) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21988))))  severity failure;
	assert RAM(21989) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21989))))  severity failure;
	assert RAM(21990) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(21990))))  severity failure;
	assert RAM(21991) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21991))))  severity failure;
	assert RAM(21992) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21992))))  severity failure;
	assert RAM(21993) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21993))))  severity failure;
	assert RAM(21994) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21994))))  severity failure;
	assert RAM(21995) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(21995))))  severity failure;
	assert RAM(21996) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21996))))  severity failure;
	assert RAM(21997) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21997))))  severity failure;
	assert RAM(21998) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21998))))  severity failure;
	assert RAM(21999) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(21999))))  severity failure;
	assert RAM(22000) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22000))))  severity failure;
	assert RAM(22001) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22001))))  severity failure;
	assert RAM(22002) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22002))))  severity failure;
	assert RAM(22003) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22003))))  severity failure;
	assert RAM(22004) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22004))))  severity failure;
	assert RAM(22005) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22005))))  severity failure;
	assert RAM(22006) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22006))))  severity failure;
	assert RAM(22007) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22007))))  severity failure;
	assert RAM(22008) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22008))))  severity failure;
	assert RAM(22009) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22009))))  severity failure;
	assert RAM(22010) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22010))))  severity failure;
	assert RAM(22011) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22011))))  severity failure;
	assert RAM(22012) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22012))))  severity failure;
	assert RAM(22013) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22013))))  severity failure;
	assert RAM(22014) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22014))))  severity failure;
	assert RAM(22015) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22015))))  severity failure;
	assert RAM(22016) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22016))))  severity failure;
	assert RAM(22017) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22017))))  severity failure;
	assert RAM(22018) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22018))))  severity failure;
	assert RAM(22019) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22019))))  severity failure;
	assert RAM(22020) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22020))))  severity failure;
	assert RAM(22021) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22021))))  severity failure;
	assert RAM(22022) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22022))))  severity failure;
	assert RAM(22023) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22023))))  severity failure;
	assert RAM(22024) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22024))))  severity failure;
	assert RAM(22025) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22025))))  severity failure;
	assert RAM(22026) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22026))))  severity failure;
	assert RAM(22027) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22027))))  severity failure;
	assert RAM(22028) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22028))))  severity failure;
	assert RAM(22029) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(22029))))  severity failure;
	assert RAM(22030) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22030))))  severity failure;
	assert RAM(22031) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(22031))))  severity failure;
	assert RAM(22032) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22032))))  severity failure;
	assert RAM(22033) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(22033))))  severity failure;
	assert RAM(22034) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22034))))  severity failure;
	assert RAM(22035) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22035))))  severity failure;
	assert RAM(22036) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22036))))  severity failure;
	assert RAM(22037) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22037))))  severity failure;
	assert RAM(22038) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22038))))  severity failure;
	assert RAM(22039) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22039))))  severity failure;
	assert RAM(22040) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22040))))  severity failure;
	assert RAM(22041) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22041))))  severity failure;
	assert RAM(22042) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22042))))  severity failure;
	assert RAM(22043) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22043))))  severity failure;
	assert RAM(22044) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(22044))))  severity failure;
	assert RAM(22045) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22045))))  severity failure;
	assert RAM(22046) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22046))))  severity failure;
	assert RAM(22047) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22047))))  severity failure;
	assert RAM(22048) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22048))))  severity failure;
	assert RAM(22049) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22049))))  severity failure;
	assert RAM(22050) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22050))))  severity failure;
	assert RAM(22051) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22051))))  severity failure;
	assert RAM(22052) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22052))))  severity failure;
	assert RAM(22053) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22053))))  severity failure;
	assert RAM(22054) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22054))))  severity failure;
	assert RAM(22055) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22055))))  severity failure;
	assert RAM(22056) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22056))))  severity failure;
	assert RAM(22057) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22057))))  severity failure;
	assert RAM(22058) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22058))))  severity failure;
	assert RAM(22059) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22059))))  severity failure;
	assert RAM(22060) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22060))))  severity failure;
	assert RAM(22061) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22061))))  severity failure;
	assert RAM(22062) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22062))))  severity failure;
	assert RAM(22063) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22063))))  severity failure;
	assert RAM(22064) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(22064))))  severity failure;
	assert RAM(22065) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22065))))  severity failure;
	assert RAM(22066) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22066))))  severity failure;
	assert RAM(22067) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22067))))  severity failure;
	assert RAM(22068) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22068))))  severity failure;
	assert RAM(22069) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22069))))  severity failure;
	assert RAM(22070) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22070))))  severity failure;
	assert RAM(22071) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22071))))  severity failure;
	assert RAM(22072) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22072))))  severity failure;
	assert RAM(22073) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22073))))  severity failure;
	assert RAM(22074) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22074))))  severity failure;
	assert RAM(22075) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22075))))  severity failure;
	assert RAM(22076) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22076))))  severity failure;
	assert RAM(22077) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22077))))  severity failure;
	assert RAM(22078) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(22078))))  severity failure;
	assert RAM(22079) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22079))))  severity failure;
	assert RAM(22080) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22080))))  severity failure;
	assert RAM(22081) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22081))))  severity failure;
	assert RAM(22082) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22082))))  severity failure;
	assert RAM(22083) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22083))))  severity failure;
	assert RAM(22084) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22084))))  severity failure;
	assert RAM(22085) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22085))))  severity failure;
	assert RAM(22086) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22086))))  severity failure;
	assert RAM(22087) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22087))))  severity failure;
	assert RAM(22088) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(22088))))  severity failure;
	assert RAM(22089) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22089))))  severity failure;
	assert RAM(22090) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22090))))  severity failure;
	assert RAM(22091) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22091))))  severity failure;
	assert RAM(22092) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22092))))  severity failure;
	assert RAM(22093) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(22093))))  severity failure;
	assert RAM(22094) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22094))))  severity failure;
	assert RAM(22095) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22095))))  severity failure;
	assert RAM(22096) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22096))))  severity failure;
	assert RAM(22097) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(22097))))  severity failure;
	assert RAM(22098) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22098))))  severity failure;
	assert RAM(22099) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(22099))))  severity failure;
	assert RAM(22100) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22100))))  severity failure;
	assert RAM(22101) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22101))))  severity failure;
	assert RAM(22102) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22102))))  severity failure;
	assert RAM(22103) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22103))))  severity failure;
	assert RAM(22104) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22104))))  severity failure;
	assert RAM(22105) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22105))))  severity failure;
	assert RAM(22106) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22106))))  severity failure;
	assert RAM(22107) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22107))))  severity failure;
	assert RAM(22108) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(22108))))  severity failure;
	assert RAM(22109) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22109))))  severity failure;
	assert RAM(22110) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(22110))))  severity failure;
	assert RAM(22111) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(22111))))  severity failure;
	assert RAM(22112) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(22112))))  severity failure;
	assert RAM(22113) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22113))))  severity failure;
	assert RAM(22114) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22114))))  severity failure;
	assert RAM(22115) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22115))))  severity failure;
	assert RAM(22116) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22116))))  severity failure;
	assert RAM(22117) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(22117))))  severity failure;
	assert RAM(22118) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22118))))  severity failure;
	assert RAM(22119) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22119))))  severity failure;
	assert RAM(22120) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22120))))  severity failure;
	assert RAM(22121) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22121))))  severity failure;
	assert RAM(22122) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22122))))  severity failure;
	assert RAM(22123) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22123))))  severity failure;
	assert RAM(22124) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(22124))))  severity failure;
	assert RAM(22125) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22125))))  severity failure;
	assert RAM(22126) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22126))))  severity failure;
	assert RAM(22127) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22127))))  severity failure;
	assert RAM(22128) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22128))))  severity failure;
	assert RAM(22129) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22129))))  severity failure;
	assert RAM(22130) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22130))))  severity failure;
	assert RAM(22131) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22131))))  severity failure;
	assert RAM(22132) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22132))))  severity failure;
	assert RAM(22133) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22133))))  severity failure;
	assert RAM(22134) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22134))))  severity failure;
	assert RAM(22135) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22135))))  severity failure;
	assert RAM(22136) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22136))))  severity failure;
	assert RAM(22137) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22137))))  severity failure;
	assert RAM(22138) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22138))))  severity failure;
	assert RAM(22139) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22139))))  severity failure;
	assert RAM(22140) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22140))))  severity failure;
	assert RAM(22141) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22141))))  severity failure;
	assert RAM(22142) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22142))))  severity failure;
	assert RAM(22143) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22143))))  severity failure;
	assert RAM(22144) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22144))))  severity failure;
	assert RAM(22145) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22145))))  severity failure;
	assert RAM(22146) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22146))))  severity failure;
	assert RAM(22147) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22147))))  severity failure;
	assert RAM(22148) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22148))))  severity failure;
	assert RAM(22149) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22149))))  severity failure;
	assert RAM(22150) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22150))))  severity failure;
	assert RAM(22151) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(22151))))  severity failure;
	assert RAM(22152) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22152))))  severity failure;
	assert RAM(22153) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22153))))  severity failure;
	assert RAM(22154) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(22154))))  severity failure;
	assert RAM(22155) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22155))))  severity failure;
	assert RAM(22156) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22156))))  severity failure;
	assert RAM(22157) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22157))))  severity failure;
	assert RAM(22158) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22158))))  severity failure;
	assert RAM(22159) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22159))))  severity failure;
	assert RAM(22160) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22160))))  severity failure;
	assert RAM(22161) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22161))))  severity failure;
	assert RAM(22162) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22162))))  severity failure;
	assert RAM(22163) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22163))))  severity failure;
	assert RAM(22164) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22164))))  severity failure;
	assert RAM(22165) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(22165))))  severity failure;
	assert RAM(22166) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22166))))  severity failure;
	assert RAM(22167) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22167))))  severity failure;
	assert RAM(22168) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22168))))  severity failure;
	assert RAM(22169) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22169))))  severity failure;
	assert RAM(22170) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22170))))  severity failure;
	assert RAM(22171) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22171))))  severity failure;
	assert RAM(22172) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22172))))  severity failure;
	assert RAM(22173) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22173))))  severity failure;
	assert RAM(22174) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22174))))  severity failure;
	assert RAM(22175) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22175))))  severity failure;
	assert RAM(22176) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22176))))  severity failure;
	assert RAM(22177) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22177))))  severity failure;
	assert RAM(22178) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22178))))  severity failure;
	assert RAM(22179) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22179))))  severity failure;
	assert RAM(22180) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(22180))))  severity failure;
	assert RAM(22181) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22181))))  severity failure;
	assert RAM(22182) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22182))))  severity failure;
	assert RAM(22183) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22183))))  severity failure;
	assert RAM(22184) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22184))))  severity failure;
	assert RAM(22185) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22185))))  severity failure;
	assert RAM(22186) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22186))))  severity failure;
	assert RAM(22187) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22187))))  severity failure;
	assert RAM(22188) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22188))))  severity failure;
	assert RAM(22189) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(22189))))  severity failure;
	assert RAM(22190) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22190))))  severity failure;
	assert RAM(22191) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22191))))  severity failure;
	assert RAM(22192) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22192))))  severity failure;
	assert RAM(22193) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(22193))))  severity failure;
	assert RAM(22194) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22194))))  severity failure;
	assert RAM(22195) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22195))))  severity failure;
	assert RAM(22196) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22196))))  severity failure;
	assert RAM(22197) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22197))))  severity failure;
	assert RAM(22198) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22198))))  severity failure;
	assert RAM(22199) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22199))))  severity failure;
	assert RAM(22200) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22200))))  severity failure;
	assert RAM(22201) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22201))))  severity failure;
	assert RAM(22202) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(22202))))  severity failure;
	assert RAM(22203) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22203))))  severity failure;
	assert RAM(22204) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(22204))))  severity failure;
	assert RAM(22205) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22205))))  severity failure;
	assert RAM(22206) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22206))))  severity failure;
	assert RAM(22207) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(22207))))  severity failure;
	assert RAM(22208) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22208))))  severity failure;
	assert RAM(22209) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22209))))  severity failure;
	assert RAM(22210) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(22210))))  severity failure;
	assert RAM(22211) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22211))))  severity failure;
	assert RAM(22212) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(22212))))  severity failure;
	assert RAM(22213) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22213))))  severity failure;
	assert RAM(22214) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22214))))  severity failure;
	assert RAM(22215) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22215))))  severity failure;
	assert RAM(22216) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(22216))))  severity failure;
	assert RAM(22217) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22217))))  severity failure;
	assert RAM(22218) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22218))))  severity failure;
	assert RAM(22219) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22219))))  severity failure;
	assert RAM(22220) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22220))))  severity failure;
	assert RAM(22221) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22221))))  severity failure;
	assert RAM(22222) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(22222))))  severity failure;
	assert RAM(22223) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22223))))  severity failure;
	assert RAM(22224) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22224))))  severity failure;
	assert RAM(22225) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22225))))  severity failure;
	assert RAM(22226) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22226))))  severity failure;
	assert RAM(22227) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22227))))  severity failure;
	assert RAM(22228) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(22228))))  severity failure;
	assert RAM(22229) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22229))))  severity failure;
	assert RAM(22230) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22230))))  severity failure;
	assert RAM(22231) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22231))))  severity failure;
	assert RAM(22232) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(22232))))  severity failure;
	assert RAM(22233) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22233))))  severity failure;
	assert RAM(22234) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22234))))  severity failure;
	assert RAM(22235) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22235))))  severity failure;
	assert RAM(22236) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22236))))  severity failure;
	assert RAM(22237) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22237))))  severity failure;
	assert RAM(22238) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22238))))  severity failure;
	assert RAM(22239) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22239))))  severity failure;
	assert RAM(22240) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22240))))  severity failure;
	assert RAM(22241) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22241))))  severity failure;
	assert RAM(22242) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22242))))  severity failure;
	assert RAM(22243) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22243))))  severity failure;
	assert RAM(22244) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22244))))  severity failure;
	assert RAM(22245) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22245))))  severity failure;
	assert RAM(22246) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22246))))  severity failure;
	assert RAM(22247) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22247))))  severity failure;
	assert RAM(22248) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22248))))  severity failure;
	assert RAM(22249) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22249))))  severity failure;
	assert RAM(22250) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22250))))  severity failure;
	assert RAM(22251) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22251))))  severity failure;
	assert RAM(22252) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22252))))  severity failure;
	assert RAM(22253) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22253))))  severity failure;
	assert RAM(22254) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22254))))  severity failure;
	assert RAM(22255) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22255))))  severity failure;
	assert RAM(22256) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22256))))  severity failure;
	assert RAM(22257) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22257))))  severity failure;
	assert RAM(22258) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22258))))  severity failure;
	assert RAM(22259) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(22259))))  severity failure;
	assert RAM(22260) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22260))))  severity failure;
	assert RAM(22261) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22261))))  severity failure;
	assert RAM(22262) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22262))))  severity failure;
	assert RAM(22263) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22263))))  severity failure;
	assert RAM(22264) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22264))))  severity failure;
	assert RAM(22265) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22265))))  severity failure;
	assert RAM(22266) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22266))))  severity failure;
	assert RAM(22267) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22267))))  severity failure;
	assert RAM(22268) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22268))))  severity failure;
	assert RAM(22269) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22269))))  severity failure;
	assert RAM(22270) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22270))))  severity failure;
	assert RAM(22271) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22271))))  severity failure;
	assert RAM(22272) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22272))))  severity failure;
	assert RAM(22273) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22273))))  severity failure;
	assert RAM(22274) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22274))))  severity failure;
	assert RAM(22275) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22275))))  severity failure;
	assert RAM(22276) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22276))))  severity failure;
	assert RAM(22277) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22277))))  severity failure;
	assert RAM(22278) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22278))))  severity failure;
	assert RAM(22279) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22279))))  severity failure;
	assert RAM(22280) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(22280))))  severity failure;
	assert RAM(22281) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(22281))))  severity failure;
	assert RAM(22282) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22282))))  severity failure;
	assert RAM(22283) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22283))))  severity failure;
	assert RAM(22284) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22284))))  severity failure;
	assert RAM(22285) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22285))))  severity failure;
	assert RAM(22286) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22286))))  severity failure;
	assert RAM(22287) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22287))))  severity failure;
	assert RAM(22288) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22288))))  severity failure;
	assert RAM(22289) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22289))))  severity failure;
	assert RAM(22290) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22290))))  severity failure;
	assert RAM(22291) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22291))))  severity failure;
	assert RAM(22292) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22292))))  severity failure;
	assert RAM(22293) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22293))))  severity failure;
	assert RAM(22294) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(22294))))  severity failure;
	assert RAM(22295) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22295))))  severity failure;
	assert RAM(22296) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22296))))  severity failure;
	assert RAM(22297) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22297))))  severity failure;
	assert RAM(22298) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22298))))  severity failure;
	assert RAM(22299) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22299))))  severity failure;
	assert RAM(22300) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22300))))  severity failure;
	assert RAM(22301) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22301))))  severity failure;
	assert RAM(22302) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22302))))  severity failure;
	assert RAM(22303) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22303))))  severity failure;
	assert RAM(22304) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22304))))  severity failure;
	assert RAM(22305) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22305))))  severity failure;
	assert RAM(22306) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22306))))  severity failure;
	assert RAM(22307) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22307))))  severity failure;
	assert RAM(22308) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22308))))  severity failure;
	assert RAM(22309) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22309))))  severity failure;
	assert RAM(22310) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22310))))  severity failure;
	assert RAM(22311) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22311))))  severity failure;
	assert RAM(22312) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22312))))  severity failure;
	assert RAM(22313) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22313))))  severity failure;
	assert RAM(22314) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22314))))  severity failure;
	assert RAM(22315) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22315))))  severity failure;
	assert RAM(22316) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22316))))  severity failure;
	assert RAM(22317) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22317))))  severity failure;
	assert RAM(22318) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22318))))  severity failure;
	assert RAM(22319) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22319))))  severity failure;
	assert RAM(22320) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22320))))  severity failure;
	assert RAM(22321) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(22321))))  severity failure;
	assert RAM(22322) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22322))))  severity failure;
	assert RAM(22323) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22323))))  severity failure;
	assert RAM(22324) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(22324))))  severity failure;
	assert RAM(22325) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22325))))  severity failure;
	assert RAM(22326) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22326))))  severity failure;
	assert RAM(22327) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22327))))  severity failure;
	assert RAM(22328) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22328))))  severity failure;
	assert RAM(22329) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22329))))  severity failure;
	assert RAM(22330) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22330))))  severity failure;
	assert RAM(22331) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22331))))  severity failure;
	assert RAM(22332) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(22332))))  severity failure;
	assert RAM(22333) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22333))))  severity failure;
	assert RAM(22334) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22334))))  severity failure;
	assert RAM(22335) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22335))))  severity failure;
	assert RAM(22336) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22336))))  severity failure;
	assert RAM(22337) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22337))))  severity failure;
	assert RAM(22338) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22338))))  severity failure;
	assert RAM(22339) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22339))))  severity failure;
	assert RAM(22340) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22340))))  severity failure;
	assert RAM(22341) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22341))))  severity failure;
	assert RAM(22342) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22342))))  severity failure;
	assert RAM(22343) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22343))))  severity failure;
	assert RAM(22344) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22344))))  severity failure;
	assert RAM(22345) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22345))))  severity failure;
	assert RAM(22346) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(22346))))  severity failure;
	assert RAM(22347) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22347))))  severity failure;
	assert RAM(22348) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22348))))  severity failure;
	assert RAM(22349) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22349))))  severity failure;
	assert RAM(22350) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22350))))  severity failure;
	assert RAM(22351) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22351))))  severity failure;
	assert RAM(22352) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22352))))  severity failure;
	assert RAM(22353) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22353))))  severity failure;
	assert RAM(22354) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22354))))  severity failure;
	assert RAM(22355) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22355))))  severity failure;
	assert RAM(22356) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22356))))  severity failure;
	assert RAM(22357) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22357))))  severity failure;
	assert RAM(22358) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22358))))  severity failure;
	assert RAM(22359) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22359))))  severity failure;
	assert RAM(22360) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22360))))  severity failure;
	assert RAM(22361) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22361))))  severity failure;
	assert RAM(22362) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22362))))  severity failure;
	assert RAM(22363) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22363))))  severity failure;
	assert RAM(22364) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22364))))  severity failure;
	assert RAM(22365) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22365))))  severity failure;
	assert RAM(22366) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22366))))  severity failure;
	assert RAM(22367) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22367))))  severity failure;
	assert RAM(22368) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22368))))  severity failure;
	assert RAM(22369) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22369))))  severity failure;
	assert RAM(22370) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22370))))  severity failure;
	assert RAM(22371) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22371))))  severity failure;
	assert RAM(22372) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22372))))  severity failure;
	assert RAM(22373) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22373))))  severity failure;
	assert RAM(22374) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22374))))  severity failure;
	assert RAM(22375) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22375))))  severity failure;
	assert RAM(22376) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(22376))))  severity failure;
	assert RAM(22377) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22377))))  severity failure;
	assert RAM(22378) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22378))))  severity failure;
	assert RAM(22379) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22379))))  severity failure;
	assert RAM(22380) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22380))))  severity failure;
	assert RAM(22381) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(22381))))  severity failure;
	assert RAM(22382) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22382))))  severity failure;
	assert RAM(22383) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22383))))  severity failure;
	assert RAM(22384) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22384))))  severity failure;
	assert RAM(22385) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22385))))  severity failure;
	assert RAM(22386) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22386))))  severity failure;
	assert RAM(22387) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22387))))  severity failure;
	assert RAM(22388) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22388))))  severity failure;
	assert RAM(22389) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22389))))  severity failure;
	assert RAM(22390) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22390))))  severity failure;
	assert RAM(22391) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22391))))  severity failure;
	assert RAM(22392) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22392))))  severity failure;
	assert RAM(22393) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22393))))  severity failure;
	assert RAM(22394) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(22394))))  severity failure;
	assert RAM(22395) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22395))))  severity failure;
	assert RAM(22396) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22396))))  severity failure;
	assert RAM(22397) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(22397))))  severity failure;
	assert RAM(22398) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22398))))  severity failure;
	assert RAM(22399) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22399))))  severity failure;
	assert RAM(22400) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22400))))  severity failure;
	assert RAM(22401) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22401))))  severity failure;
	assert RAM(22402) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22402))))  severity failure;
	assert RAM(22403) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(22403))))  severity failure;
	assert RAM(22404) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22404))))  severity failure;
	assert RAM(22405) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22405))))  severity failure;
	assert RAM(22406) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(22406))))  severity failure;
	assert RAM(22407) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22407))))  severity failure;
	assert RAM(22408) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22408))))  severity failure;
	assert RAM(22409) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22409))))  severity failure;
	assert RAM(22410) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22410))))  severity failure;
	assert RAM(22411) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22411))))  severity failure;
	assert RAM(22412) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(22412))))  severity failure;
	assert RAM(22413) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22413))))  severity failure;
	assert RAM(22414) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(22414))))  severity failure;
	assert RAM(22415) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22415))))  severity failure;
	assert RAM(22416) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(22416))))  severity failure;
	assert RAM(22417) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(22417))))  severity failure;
	assert RAM(22418) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22418))))  severity failure;
	assert RAM(22419) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22419))))  severity failure;
	assert RAM(22420) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22420))))  severity failure;
	assert RAM(22421) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22421))))  severity failure;
	assert RAM(22422) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(22422))))  severity failure;
	assert RAM(22423) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22423))))  severity failure;
	assert RAM(22424) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22424))))  severity failure;
	assert RAM(22425) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22425))))  severity failure;
	assert RAM(22426) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22426))))  severity failure;
	assert RAM(22427) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22427))))  severity failure;
	assert RAM(22428) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22428))))  severity failure;
	assert RAM(22429) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22429))))  severity failure;
	assert RAM(22430) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22430))))  severity failure;
	assert RAM(22431) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22431))))  severity failure;
	assert RAM(22432) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(22432))))  severity failure;
	assert RAM(22433) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22433))))  severity failure;
	assert RAM(22434) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22434))))  severity failure;
	assert RAM(22435) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22435))))  severity failure;
	assert RAM(22436) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22436))))  severity failure;
	assert RAM(22437) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22437))))  severity failure;
	assert RAM(22438) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22438))))  severity failure;
	assert RAM(22439) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22439))))  severity failure;
	assert RAM(22440) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(22440))))  severity failure;
	assert RAM(22441) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22441))))  severity failure;
	assert RAM(22442) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22442))))  severity failure;
	assert RAM(22443) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22443))))  severity failure;
	assert RAM(22444) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22444))))  severity failure;
	assert RAM(22445) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22445))))  severity failure;
	assert RAM(22446) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22446))))  severity failure;
	assert RAM(22447) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22447))))  severity failure;
	assert RAM(22448) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(22448))))  severity failure;
	assert RAM(22449) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22449))))  severity failure;
	assert RAM(22450) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22450))))  severity failure;
	assert RAM(22451) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22451))))  severity failure;
	assert RAM(22452) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22452))))  severity failure;
	assert RAM(22453) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22453))))  severity failure;
	assert RAM(22454) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22454))))  severity failure;
	assert RAM(22455) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22455))))  severity failure;
	assert RAM(22456) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22456))))  severity failure;
	assert RAM(22457) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22457))))  severity failure;
	assert RAM(22458) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22458))))  severity failure;
	assert RAM(22459) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22459))))  severity failure;
	assert RAM(22460) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22460))))  severity failure;
	assert RAM(22461) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22461))))  severity failure;
	assert RAM(22462) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22462))))  severity failure;
	assert RAM(22463) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22463))))  severity failure;
	assert RAM(22464) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(22464))))  severity failure;
	assert RAM(22465) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22465))))  severity failure;
	assert RAM(22466) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22466))))  severity failure;
	assert RAM(22467) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22467))))  severity failure;
	assert RAM(22468) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22468))))  severity failure;
	assert RAM(22469) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22469))))  severity failure;
	assert RAM(22470) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22470))))  severity failure;
	assert RAM(22471) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22471))))  severity failure;
	assert RAM(22472) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(22472))))  severity failure;
	assert RAM(22473) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22473))))  severity failure;
	assert RAM(22474) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22474))))  severity failure;
	assert RAM(22475) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22475))))  severity failure;
	assert RAM(22476) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22476))))  severity failure;
	assert RAM(22477) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22477))))  severity failure;
	assert RAM(22478) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22478))))  severity failure;
	assert RAM(22479) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22479))))  severity failure;
	assert RAM(22480) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22480))))  severity failure;
	assert RAM(22481) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22481))))  severity failure;
	assert RAM(22482) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22482))))  severity failure;
	assert RAM(22483) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22483))))  severity failure;
	assert RAM(22484) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22484))))  severity failure;
	assert RAM(22485) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(22485))))  severity failure;
	assert RAM(22486) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22486))))  severity failure;
	assert RAM(22487) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22487))))  severity failure;
	assert RAM(22488) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22488))))  severity failure;
	assert RAM(22489) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22489))))  severity failure;
	assert RAM(22490) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22490))))  severity failure;
	assert RAM(22491) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22491))))  severity failure;
	assert RAM(22492) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22492))))  severity failure;
	assert RAM(22493) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22493))))  severity failure;
	assert RAM(22494) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(22494))))  severity failure;
	assert RAM(22495) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22495))))  severity failure;
	assert RAM(22496) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22496))))  severity failure;
	assert RAM(22497) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(22497))))  severity failure;
	assert RAM(22498) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(22498))))  severity failure;
	assert RAM(22499) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22499))))  severity failure;
	assert RAM(22500) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22500))))  severity failure;
	assert RAM(22501) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22501))))  severity failure;
	assert RAM(22502) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22502))))  severity failure;
	assert RAM(22503) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22503))))  severity failure;
	assert RAM(22504) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22504))))  severity failure;
	assert RAM(22505) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22505))))  severity failure;
	assert RAM(22506) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22506))))  severity failure;
	assert RAM(22507) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22507))))  severity failure;
	assert RAM(22508) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22508))))  severity failure;
	assert RAM(22509) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22509))))  severity failure;
	assert RAM(22510) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22510))))  severity failure;
	assert RAM(22511) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22511))))  severity failure;
	assert RAM(22512) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(22512))))  severity failure;
	assert RAM(22513) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22513))))  severity failure;
	assert RAM(22514) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22514))))  severity failure;
	assert RAM(22515) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22515))))  severity failure;
	assert RAM(22516) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22516))))  severity failure;
	assert RAM(22517) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22517))))  severity failure;
	assert RAM(22518) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(22518))))  severity failure;
	assert RAM(22519) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22519))))  severity failure;
	assert RAM(22520) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22520))))  severity failure;
	assert RAM(22521) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(22521))))  severity failure;
	assert RAM(22522) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(22522))))  severity failure;
	assert RAM(22523) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22523))))  severity failure;
	assert RAM(22524) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22524))))  severity failure;
	assert RAM(22525) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22525))))  severity failure;
	assert RAM(22526) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22526))))  severity failure;
	assert RAM(22527) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22527))))  severity failure;
	assert RAM(22528) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22528))))  severity failure;
	assert RAM(22529) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22529))))  severity failure;
	assert RAM(22530) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22530))))  severity failure;
	assert RAM(22531) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22531))))  severity failure;
	assert RAM(22532) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22532))))  severity failure;
	assert RAM(22533) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22533))))  severity failure;
	assert RAM(22534) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22534))))  severity failure;
	assert RAM(22535) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22535))))  severity failure;
	assert RAM(22536) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22536))))  severity failure;
	assert RAM(22537) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22537))))  severity failure;
	assert RAM(22538) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22538))))  severity failure;
	assert RAM(22539) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(22539))))  severity failure;
	assert RAM(22540) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22540))))  severity failure;
	assert RAM(22541) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22541))))  severity failure;
	assert RAM(22542) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22542))))  severity failure;
	assert RAM(22543) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(22543))))  severity failure;
	assert RAM(22544) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22544))))  severity failure;
	assert RAM(22545) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22545))))  severity failure;
	assert RAM(22546) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22546))))  severity failure;
	assert RAM(22547) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22547))))  severity failure;
	assert RAM(22548) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22548))))  severity failure;
	assert RAM(22549) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22549))))  severity failure;
	assert RAM(22550) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(22550))))  severity failure;
	assert RAM(22551) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22551))))  severity failure;
	assert RAM(22552) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22552))))  severity failure;
	assert RAM(22553) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22553))))  severity failure;
	assert RAM(22554) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22554))))  severity failure;
	assert RAM(22555) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22555))))  severity failure;
	assert RAM(22556) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22556))))  severity failure;
	assert RAM(22557) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22557))))  severity failure;
	assert RAM(22558) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22558))))  severity failure;
	assert RAM(22559) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(22559))))  severity failure;
	assert RAM(22560) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22560))))  severity failure;
	assert RAM(22561) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22561))))  severity failure;
	assert RAM(22562) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22562))))  severity failure;
	assert RAM(22563) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22563))))  severity failure;
	assert RAM(22564) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22564))))  severity failure;
	assert RAM(22565) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22565))))  severity failure;
	assert RAM(22566) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22566))))  severity failure;
	assert RAM(22567) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22567))))  severity failure;
	assert RAM(22568) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22568))))  severity failure;
	assert RAM(22569) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22569))))  severity failure;
	assert RAM(22570) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22570))))  severity failure;
	assert RAM(22571) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22571))))  severity failure;
	assert RAM(22572) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22572))))  severity failure;
	assert RAM(22573) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22573))))  severity failure;
	assert RAM(22574) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22574))))  severity failure;
	assert RAM(22575) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22575))))  severity failure;
	assert RAM(22576) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22576))))  severity failure;
	assert RAM(22577) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22577))))  severity failure;
	assert RAM(22578) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22578))))  severity failure;
	assert RAM(22579) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22579))))  severity failure;
	assert RAM(22580) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22580))))  severity failure;
	assert RAM(22581) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22581))))  severity failure;
	assert RAM(22582) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22582))))  severity failure;
	assert RAM(22583) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22583))))  severity failure;
	assert RAM(22584) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22584))))  severity failure;
	assert RAM(22585) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(22585))))  severity failure;
	assert RAM(22586) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22586))))  severity failure;
	assert RAM(22587) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22587))))  severity failure;
	assert RAM(22588) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22588))))  severity failure;
	assert RAM(22589) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22589))))  severity failure;
	assert RAM(22590) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22590))))  severity failure;
	assert RAM(22591) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(22591))))  severity failure;
	assert RAM(22592) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22592))))  severity failure;
	assert RAM(22593) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22593))))  severity failure;
	assert RAM(22594) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22594))))  severity failure;
	assert RAM(22595) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22595))))  severity failure;
	assert RAM(22596) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22596))))  severity failure;
	assert RAM(22597) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22597))))  severity failure;
	assert RAM(22598) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22598))))  severity failure;
	assert RAM(22599) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22599))))  severity failure;
	assert RAM(22600) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22600))))  severity failure;
	assert RAM(22601) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22601))))  severity failure;
	assert RAM(22602) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22602))))  severity failure;
	assert RAM(22603) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(22603))))  severity failure;
	assert RAM(22604) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22604))))  severity failure;
	assert RAM(22605) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22605))))  severity failure;
	assert RAM(22606) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22606))))  severity failure;
	assert RAM(22607) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22607))))  severity failure;
	assert RAM(22608) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22608))))  severity failure;
	assert RAM(22609) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22609))))  severity failure;
	assert RAM(22610) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22610))))  severity failure;
	assert RAM(22611) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22611))))  severity failure;
	assert RAM(22612) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(22612))))  severity failure;
	assert RAM(22613) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22613))))  severity failure;
	assert RAM(22614) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22614))))  severity failure;
	assert RAM(22615) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22615))))  severity failure;
	assert RAM(22616) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22616))))  severity failure;
	assert RAM(22617) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22617))))  severity failure;
	assert RAM(22618) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22618))))  severity failure;
	assert RAM(22619) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22619))))  severity failure;
	assert RAM(22620) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22620))))  severity failure;
	assert RAM(22621) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22621))))  severity failure;
	assert RAM(22622) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22622))))  severity failure;
	assert RAM(22623) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22623))))  severity failure;
	assert RAM(22624) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22624))))  severity failure;
	assert RAM(22625) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22625))))  severity failure;
	assert RAM(22626) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(22626))))  severity failure;
	assert RAM(22627) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22627))))  severity failure;
	assert RAM(22628) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22628))))  severity failure;
	assert RAM(22629) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(22629))))  severity failure;
	assert RAM(22630) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22630))))  severity failure;
	assert RAM(22631) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22631))))  severity failure;
	assert RAM(22632) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22632))))  severity failure;
	assert RAM(22633) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22633))))  severity failure;
	assert RAM(22634) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(22634))))  severity failure;
	assert RAM(22635) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22635))))  severity failure;
	assert RAM(22636) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22636))))  severity failure;
	assert RAM(22637) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22637))))  severity failure;
	assert RAM(22638) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22638))))  severity failure;
	assert RAM(22639) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(22639))))  severity failure;
	assert RAM(22640) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(22640))))  severity failure;
	assert RAM(22641) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22641))))  severity failure;
	assert RAM(22642) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22642))))  severity failure;
	assert RAM(22643) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22643))))  severity failure;
	assert RAM(22644) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22644))))  severity failure;
	assert RAM(22645) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22645))))  severity failure;
	assert RAM(22646) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22646))))  severity failure;
	assert RAM(22647) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22647))))  severity failure;
	assert RAM(22648) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22648))))  severity failure;
	assert RAM(22649) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22649))))  severity failure;
	assert RAM(22650) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22650))))  severity failure;
	assert RAM(22651) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22651))))  severity failure;
	assert RAM(22652) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(22652))))  severity failure;
	assert RAM(22653) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22653))))  severity failure;
	assert RAM(22654) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22654))))  severity failure;
	assert RAM(22655) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22655))))  severity failure;
	assert RAM(22656) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(22656))))  severity failure;
	assert RAM(22657) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22657))))  severity failure;
	assert RAM(22658) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22658))))  severity failure;
	assert RAM(22659) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22659))))  severity failure;
	assert RAM(22660) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22660))))  severity failure;
	assert RAM(22661) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22661))))  severity failure;
	assert RAM(22662) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22662))))  severity failure;
	assert RAM(22663) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22663))))  severity failure;
	assert RAM(22664) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22664))))  severity failure;
	assert RAM(22665) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22665))))  severity failure;
	assert RAM(22666) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22666))))  severity failure;
	assert RAM(22667) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22667))))  severity failure;
	assert RAM(22668) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22668))))  severity failure;
	assert RAM(22669) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22669))))  severity failure;
	assert RAM(22670) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22670))))  severity failure;
	assert RAM(22671) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22671))))  severity failure;
	assert RAM(22672) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22672))))  severity failure;
	assert RAM(22673) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22673))))  severity failure;
	assert RAM(22674) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22674))))  severity failure;
	assert RAM(22675) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22675))))  severity failure;
	assert RAM(22676) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(22676))))  severity failure;
	assert RAM(22677) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22677))))  severity failure;
	assert RAM(22678) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22678))))  severity failure;
	assert RAM(22679) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(22679))))  severity failure;
	assert RAM(22680) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22680))))  severity failure;
	assert RAM(22681) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22681))))  severity failure;
	assert RAM(22682) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22682))))  severity failure;
	assert RAM(22683) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22683))))  severity failure;
	assert RAM(22684) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22684))))  severity failure;
	assert RAM(22685) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22685))))  severity failure;
	assert RAM(22686) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22686))))  severity failure;
	assert RAM(22687) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22687))))  severity failure;
	assert RAM(22688) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22688))))  severity failure;
	assert RAM(22689) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22689))))  severity failure;
	assert RAM(22690) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(22690))))  severity failure;
	assert RAM(22691) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22691))))  severity failure;
	assert RAM(22692) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22692))))  severity failure;
	assert RAM(22693) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22693))))  severity failure;
	assert RAM(22694) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22694))))  severity failure;
	assert RAM(22695) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22695))))  severity failure;
	assert RAM(22696) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22696))))  severity failure;
	assert RAM(22697) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22697))))  severity failure;
	assert RAM(22698) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22698))))  severity failure;
	assert RAM(22699) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(22699))))  severity failure;
	assert RAM(22700) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22700))))  severity failure;
	assert RAM(22701) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22701))))  severity failure;
	assert RAM(22702) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(22702))))  severity failure;
	assert RAM(22703) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22703))))  severity failure;
	assert RAM(22704) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22704))))  severity failure;
	assert RAM(22705) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22705))))  severity failure;
	assert RAM(22706) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22706))))  severity failure;
	assert RAM(22707) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22707))))  severity failure;
	assert RAM(22708) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22708))))  severity failure;
	assert RAM(22709) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(22709))))  severity failure;
	assert RAM(22710) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(22710))))  severity failure;
	assert RAM(22711) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22711))))  severity failure;
	assert RAM(22712) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22712))))  severity failure;
	assert RAM(22713) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22713))))  severity failure;
	assert RAM(22714) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22714))))  severity failure;
	assert RAM(22715) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22715))))  severity failure;
	assert RAM(22716) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22716))))  severity failure;
	assert RAM(22717) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22717))))  severity failure;
	assert RAM(22718) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22718))))  severity failure;
	assert RAM(22719) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22719))))  severity failure;
	assert RAM(22720) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22720))))  severity failure;
	assert RAM(22721) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22721))))  severity failure;
	assert RAM(22722) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(22722))))  severity failure;
	assert RAM(22723) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22723))))  severity failure;
	assert RAM(22724) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(22724))))  severity failure;
	assert RAM(22725) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22725))))  severity failure;
	assert RAM(22726) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22726))))  severity failure;
	assert RAM(22727) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22727))))  severity failure;
	assert RAM(22728) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22728))))  severity failure;
	assert RAM(22729) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22729))))  severity failure;
	assert RAM(22730) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22730))))  severity failure;
	assert RAM(22731) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(22731))))  severity failure;
	assert RAM(22732) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22732))))  severity failure;
	assert RAM(22733) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22733))))  severity failure;
	assert RAM(22734) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22734))))  severity failure;
	assert RAM(22735) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22735))))  severity failure;
	assert RAM(22736) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22736))))  severity failure;
	assert RAM(22737) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22737))))  severity failure;
	assert RAM(22738) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22738))))  severity failure;
	assert RAM(22739) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22739))))  severity failure;
	assert RAM(22740) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22740))))  severity failure;
	assert RAM(22741) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22741))))  severity failure;
	assert RAM(22742) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22742))))  severity failure;
	assert RAM(22743) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22743))))  severity failure;
	assert RAM(22744) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22744))))  severity failure;
	assert RAM(22745) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22745))))  severity failure;
	assert RAM(22746) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22746))))  severity failure;
	assert RAM(22747) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22747))))  severity failure;
	assert RAM(22748) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22748))))  severity failure;
	assert RAM(22749) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22749))))  severity failure;
	assert RAM(22750) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22750))))  severity failure;
	assert RAM(22751) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22751))))  severity failure;
	assert RAM(22752) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22752))))  severity failure;
	assert RAM(22753) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22753))))  severity failure;
	assert RAM(22754) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22754))))  severity failure;
	assert RAM(22755) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22755))))  severity failure;
	assert RAM(22756) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22756))))  severity failure;
	assert RAM(22757) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22757))))  severity failure;
	assert RAM(22758) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22758))))  severity failure;
	assert RAM(22759) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22759))))  severity failure;
	assert RAM(22760) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22760))))  severity failure;
	assert RAM(22761) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22761))))  severity failure;
	assert RAM(22762) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22762))))  severity failure;
	assert RAM(22763) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22763))))  severity failure;
	assert RAM(22764) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22764))))  severity failure;
	assert RAM(22765) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22765))))  severity failure;
	assert RAM(22766) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22766))))  severity failure;
	assert RAM(22767) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(22767))))  severity failure;
	assert RAM(22768) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22768))))  severity failure;
	assert RAM(22769) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22769))))  severity failure;
	assert RAM(22770) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22770))))  severity failure;
	assert RAM(22771) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22771))))  severity failure;
	assert RAM(22772) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22772))))  severity failure;
	assert RAM(22773) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(22773))))  severity failure;
	assert RAM(22774) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22774))))  severity failure;
	assert RAM(22775) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22775))))  severity failure;
	assert RAM(22776) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22776))))  severity failure;
	assert RAM(22777) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22777))))  severity failure;
	assert RAM(22778) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22778))))  severity failure;
	assert RAM(22779) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22779))))  severity failure;
	assert RAM(22780) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22780))))  severity failure;
	assert RAM(22781) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22781))))  severity failure;
	assert RAM(22782) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22782))))  severity failure;
	assert RAM(22783) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22783))))  severity failure;
	assert RAM(22784) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22784))))  severity failure;
	assert RAM(22785) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22785))))  severity failure;
	assert RAM(22786) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22786))))  severity failure;
	assert RAM(22787) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22787))))  severity failure;
	assert RAM(22788) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22788))))  severity failure;
	assert RAM(22789) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22789))))  severity failure;
	assert RAM(22790) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22790))))  severity failure;
	assert RAM(22791) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22791))))  severity failure;
	assert RAM(22792) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22792))))  severity failure;
	assert RAM(22793) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22793))))  severity failure;
	assert RAM(22794) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22794))))  severity failure;
	assert RAM(22795) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22795))))  severity failure;
	assert RAM(22796) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22796))))  severity failure;
	assert RAM(22797) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(22797))))  severity failure;
	assert RAM(22798) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22798))))  severity failure;
	assert RAM(22799) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22799))))  severity failure;
	assert RAM(22800) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22800))))  severity failure;
	assert RAM(22801) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22801))))  severity failure;
	assert RAM(22802) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(22802))))  severity failure;
	assert RAM(22803) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22803))))  severity failure;
	assert RAM(22804) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22804))))  severity failure;
	assert RAM(22805) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22805))))  severity failure;
	assert RAM(22806) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22806))))  severity failure;
	assert RAM(22807) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22807))))  severity failure;
	assert RAM(22808) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22808))))  severity failure;
	assert RAM(22809) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22809))))  severity failure;
	assert RAM(22810) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22810))))  severity failure;
	assert RAM(22811) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22811))))  severity failure;
	assert RAM(22812) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22812))))  severity failure;
	assert RAM(22813) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22813))))  severity failure;
	assert RAM(22814) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22814))))  severity failure;
	assert RAM(22815) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22815))))  severity failure;
	assert RAM(22816) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22816))))  severity failure;
	assert RAM(22817) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22817))))  severity failure;
	assert RAM(22818) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22818))))  severity failure;
	assert RAM(22819) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22819))))  severity failure;
	assert RAM(22820) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(22820))))  severity failure;
	assert RAM(22821) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22821))))  severity failure;
	assert RAM(22822) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22822))))  severity failure;
	assert RAM(22823) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22823))))  severity failure;
	assert RAM(22824) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22824))))  severity failure;
	assert RAM(22825) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22825))))  severity failure;
	assert RAM(22826) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22826))))  severity failure;
	assert RAM(22827) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22827))))  severity failure;
	assert RAM(22828) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22828))))  severity failure;
	assert RAM(22829) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(22829))))  severity failure;
	assert RAM(22830) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22830))))  severity failure;
	assert RAM(22831) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(22831))))  severity failure;
	assert RAM(22832) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22832))))  severity failure;
	assert RAM(22833) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22833))))  severity failure;
	assert RAM(22834) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22834))))  severity failure;
	assert RAM(22835) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22835))))  severity failure;
	assert RAM(22836) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22836))))  severity failure;
	assert RAM(22837) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22837))))  severity failure;
	assert RAM(22838) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22838))))  severity failure;
	assert RAM(22839) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22839))))  severity failure;
	assert RAM(22840) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22840))))  severity failure;
	assert RAM(22841) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22841))))  severity failure;
	assert RAM(22842) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22842))))  severity failure;
	assert RAM(22843) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22843))))  severity failure;
	assert RAM(22844) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22844))))  severity failure;
	assert RAM(22845) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22845))))  severity failure;
	assert RAM(22846) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(22846))))  severity failure;
	assert RAM(22847) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22847))))  severity failure;
	assert RAM(22848) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22848))))  severity failure;
	assert RAM(22849) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22849))))  severity failure;
	assert RAM(22850) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22850))))  severity failure;
	assert RAM(22851) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22851))))  severity failure;
	assert RAM(22852) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22852))))  severity failure;
	assert RAM(22853) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22853))))  severity failure;
	assert RAM(22854) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22854))))  severity failure;
	assert RAM(22855) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(22855))))  severity failure;
	assert RAM(22856) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22856))))  severity failure;
	assert RAM(22857) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22857))))  severity failure;
	assert RAM(22858) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22858))))  severity failure;
	assert RAM(22859) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22859))))  severity failure;
	assert RAM(22860) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22860))))  severity failure;
	assert RAM(22861) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(22861))))  severity failure;
	assert RAM(22862) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22862))))  severity failure;
	assert RAM(22863) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22863))))  severity failure;
	assert RAM(22864) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22864))))  severity failure;
	assert RAM(22865) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(22865))))  severity failure;
	assert RAM(22866) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22866))))  severity failure;
	assert RAM(22867) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22867))))  severity failure;
	assert RAM(22868) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22868))))  severity failure;
	assert RAM(22869) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22869))))  severity failure;
	assert RAM(22870) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22870))))  severity failure;
	assert RAM(22871) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22871))))  severity failure;
	assert RAM(22872) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22872))))  severity failure;
	assert RAM(22873) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22873))))  severity failure;
	assert RAM(22874) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22874))))  severity failure;
	assert RAM(22875) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(22875))))  severity failure;
	assert RAM(22876) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(22876))))  severity failure;
	assert RAM(22877) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22877))))  severity failure;
	assert RAM(22878) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(22878))))  severity failure;
	assert RAM(22879) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(22879))))  severity failure;
	assert RAM(22880) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22880))))  severity failure;
	assert RAM(22881) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22881))))  severity failure;
	assert RAM(22882) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22882))))  severity failure;
	assert RAM(22883) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22883))))  severity failure;
	assert RAM(22884) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22884))))  severity failure;
	assert RAM(22885) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22885))))  severity failure;
	assert RAM(22886) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22886))))  severity failure;
	assert RAM(22887) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22887))))  severity failure;
	assert RAM(22888) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22888))))  severity failure;
	assert RAM(22889) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22889))))  severity failure;
	assert RAM(22890) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22890))))  severity failure;
	assert RAM(22891) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22891))))  severity failure;
	assert RAM(22892) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22892))))  severity failure;
	assert RAM(22893) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22893))))  severity failure;
	assert RAM(22894) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22894))))  severity failure;
	assert RAM(22895) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22895))))  severity failure;
	assert RAM(22896) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22896))))  severity failure;
	assert RAM(22897) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22897))))  severity failure;
	assert RAM(22898) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22898))))  severity failure;
	assert RAM(22899) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22899))))  severity failure;
	assert RAM(22900) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22900))))  severity failure;
	assert RAM(22901) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22901))))  severity failure;
	assert RAM(22902) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22902))))  severity failure;
	assert RAM(22903) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22903))))  severity failure;
	assert RAM(22904) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(22904))))  severity failure;
	assert RAM(22905) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22905))))  severity failure;
	assert RAM(22906) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22906))))  severity failure;
	assert RAM(22907) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22907))))  severity failure;
	assert RAM(22908) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22908))))  severity failure;
	assert RAM(22909) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22909))))  severity failure;
	assert RAM(22910) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22910))))  severity failure;
	assert RAM(22911) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22911))))  severity failure;
	assert RAM(22912) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22912))))  severity failure;
	assert RAM(22913) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22913))))  severity failure;
	assert RAM(22914) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22914))))  severity failure;
	assert RAM(22915) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22915))))  severity failure;
	assert RAM(22916) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(22916))))  severity failure;
	assert RAM(22917) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22917))))  severity failure;
	assert RAM(22918) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(22918))))  severity failure;
	assert RAM(22919) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22919))))  severity failure;
	assert RAM(22920) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22920))))  severity failure;
	assert RAM(22921) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22921))))  severity failure;
	assert RAM(22922) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22922))))  severity failure;
	assert RAM(22923) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22923))))  severity failure;
	assert RAM(22924) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22924))))  severity failure;
	assert RAM(22925) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22925))))  severity failure;
	assert RAM(22926) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22926))))  severity failure;
	assert RAM(22927) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(22927))))  severity failure;
	assert RAM(22928) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22928))))  severity failure;
	assert RAM(22929) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22929))))  severity failure;
	assert RAM(22930) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22930))))  severity failure;
	assert RAM(22931) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22931))))  severity failure;
	assert RAM(22932) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(22932))))  severity failure;
	assert RAM(22933) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(22933))))  severity failure;
	assert RAM(22934) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22934))))  severity failure;
	assert RAM(22935) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22935))))  severity failure;
	assert RAM(22936) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22936))))  severity failure;
	assert RAM(22937) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22937))))  severity failure;
	assert RAM(22938) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22938))))  severity failure;
	assert RAM(22939) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22939))))  severity failure;
	assert RAM(22940) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22940))))  severity failure;
	assert RAM(22941) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22941))))  severity failure;
	assert RAM(22942) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22942))))  severity failure;
	assert RAM(22943) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22943))))  severity failure;
	assert RAM(22944) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22944))))  severity failure;
	assert RAM(22945) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22945))))  severity failure;
	assert RAM(22946) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22946))))  severity failure;
	assert RAM(22947) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22947))))  severity failure;
	assert RAM(22948) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22948))))  severity failure;
	assert RAM(22949) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22949))))  severity failure;
	assert RAM(22950) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22950))))  severity failure;
	assert RAM(22951) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22951))))  severity failure;
	assert RAM(22952) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22952))))  severity failure;
	assert RAM(22953) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22953))))  severity failure;
	assert RAM(22954) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22954))))  severity failure;
	assert RAM(22955) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22955))))  severity failure;
	assert RAM(22956) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22956))))  severity failure;
	assert RAM(22957) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22957))))  severity failure;
	assert RAM(22958) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22958))))  severity failure;
	assert RAM(22959) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22959))))  severity failure;
	assert RAM(22960) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22960))))  severity failure;
	assert RAM(22961) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22961))))  severity failure;
	assert RAM(22962) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22962))))  severity failure;
	assert RAM(22963) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22963))))  severity failure;
	assert RAM(22964) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(22964))))  severity failure;
	assert RAM(22965) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22965))))  severity failure;
	assert RAM(22966) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22966))))  severity failure;
	assert RAM(22967) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22967))))  severity failure;
	assert RAM(22968) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(22968))))  severity failure;
	assert RAM(22969) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(22969))))  severity failure;
	assert RAM(22970) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22970))))  severity failure;
	assert RAM(22971) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(22971))))  severity failure;
	assert RAM(22972) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(22972))))  severity failure;
	assert RAM(22973) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22973))))  severity failure;
	assert RAM(22974) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22974))))  severity failure;
	assert RAM(22975) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22975))))  severity failure;
	assert RAM(22976) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22976))))  severity failure;
	assert RAM(22977) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22977))))  severity failure;
	assert RAM(22978) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22978))))  severity failure;
	assert RAM(22979) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22979))))  severity failure;
	assert RAM(22980) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22980))))  severity failure;
	assert RAM(22981) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22981))))  severity failure;
	assert RAM(22982) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22982))))  severity failure;
	assert RAM(22983) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22983))))  severity failure;
	assert RAM(22984) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22984))))  severity failure;
	assert RAM(22985) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22985))))  severity failure;
	assert RAM(22986) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22986))))  severity failure;
	assert RAM(22987) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22987))))  severity failure;
	assert RAM(22988) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22988))))  severity failure;
	assert RAM(22989) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22989))))  severity failure;
	assert RAM(22990) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22990))))  severity failure;
	assert RAM(22991) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22991))))  severity failure;
	assert RAM(22992) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22992))))  severity failure;
	assert RAM(22993) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22993))))  severity failure;
	assert RAM(22994) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22994))))  severity failure;
	assert RAM(22995) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22995))))  severity failure;
	assert RAM(22996) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22996))))  severity failure;
	assert RAM(22997) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22997))))  severity failure;
	assert RAM(22998) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22998))))  severity failure;
	assert RAM(22999) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22999))))  severity failure;
	assert RAM(23000) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23000))))  severity failure;
	assert RAM(23001) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(23001))))  severity failure;
	assert RAM(23002) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23002))))  severity failure;
	assert RAM(23003) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23003))))  severity failure;
	assert RAM(23004) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23004))))  severity failure;
	assert RAM(23005) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(23005))))  severity failure;
	assert RAM(23006) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23006))))  severity failure;
	assert RAM(23007) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23007))))  severity failure;
	assert RAM(23008) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(23008))))  severity failure;
	assert RAM(23009) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(23009))))  severity failure;
	assert RAM(23010) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23010))))  severity failure;
	assert RAM(23011) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(23011))))  severity failure;
	assert RAM(23012) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(23012))))  severity failure;
	assert RAM(23013) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23013))))  severity failure;
	assert RAM(23014) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(23014))))  severity failure;
	assert RAM(23015) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23015))))  severity failure;
	assert RAM(23016) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(23016))))  severity failure;
	assert RAM(23017) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(23017))))  severity failure;
	assert RAM(23018) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23018))))  severity failure;
	assert RAM(23019) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23019))))  severity failure;
	assert RAM(23020) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(23020))))  severity failure;
	assert RAM(23021) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23021))))  severity failure;
	assert RAM(23022) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(23022))))  severity failure;
	assert RAM(23023) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23023))))  severity failure;
	assert RAM(23024) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(23024))))  severity failure;
	assert RAM(23025) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(23025))))  severity failure;
	assert RAM(23026) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23026))))  severity failure;
	assert RAM(23027) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23027))))  severity failure;
	assert RAM(23028) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23028))))  severity failure;
	assert RAM(23029) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23029))))  severity failure;
	assert RAM(23030) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23030))))  severity failure;
	assert RAM(23031) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23031))))  severity failure;
	assert RAM(23032) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(23032))))  severity failure;
	assert RAM(23033) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(23033))))  severity failure;
	assert RAM(23034) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(23034))))  severity failure;
	assert RAM(23035) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23035))))  severity failure;
	assert RAM(23036) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(23036))))  severity failure;
	assert RAM(23037) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23037))))  severity failure;
	assert RAM(23038) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23038))))  severity failure;
	assert RAM(23039) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(23039))))  severity failure;
	assert RAM(23040) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23040))))  severity failure;
	assert RAM(23041) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(23041))))  severity failure;
	assert RAM(23042) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23042))))  severity failure;
	assert RAM(23043) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23043))))  severity failure;
	assert RAM(23044) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23044))))  severity failure;
	assert RAM(23045) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(23045))))  severity failure;
	assert RAM(23046) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23046))))  severity failure;
	assert RAM(23047) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23047))))  severity failure;
	assert RAM(23048) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23048))))  severity failure;
	assert RAM(23049) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23049))))  severity failure;
	assert RAM(23050) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(23050))))  severity failure;
	assert RAM(23051) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23051))))  severity failure;
	assert RAM(23052) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23052))))  severity failure;
	assert RAM(23053) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23053))))  severity failure;
	assert RAM(23054) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23054))))  severity failure;
	assert RAM(23055) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(23055))))  severity failure;
	assert RAM(23056) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23056))))  severity failure;
	assert RAM(23057) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23057))))  severity failure;
	assert RAM(23058) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23058))))  severity failure;
	assert RAM(23059) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(23059))))  severity failure;
	assert RAM(23060) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(23060))))  severity failure;
	assert RAM(23061) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23061))))  severity failure;
	assert RAM(23062) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23062))))  severity failure;
	assert RAM(23063) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(23063))))  severity failure;
	assert RAM(23064) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(23064))))  severity failure;
	assert RAM(23065) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23065))))  severity failure;
	assert RAM(23066) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23066))))  severity failure;
	assert RAM(23067) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(23067))))  severity failure;
	assert RAM(23068) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(23068))))  severity failure;
	assert RAM(23069) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(23069))))  severity failure;
	assert RAM(23070) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23070))))  severity failure;
	assert RAM(23071) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(23071))))  severity failure;
	assert RAM(23072) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23072))))  severity failure;
	assert RAM(23073) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23073))))  severity failure;
	assert RAM(23074) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(23074))))  severity failure;
	assert RAM(23075) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23075))))  severity failure;
	assert RAM(23076) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23076))))  severity failure;
	assert RAM(23077) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23077))))  severity failure;
	assert RAM(23078) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23078))))  severity failure;
	assert RAM(23079) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23079))))  severity failure;
	assert RAM(23080) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(23080))))  severity failure;
	assert RAM(23081) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23081))))  severity failure;
	assert RAM(23082) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23082))))  severity failure;
	assert RAM(23083) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23083))))  severity failure;
	assert RAM(23084) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23084))))  severity failure;
	assert RAM(23085) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(23085))))  severity failure;
	assert RAM(23086) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23086))))  severity failure;
	assert RAM(23087) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(23087))))  severity failure;
	assert RAM(23088) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(23088))))  severity failure;
	assert RAM(23089) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23089))))  severity failure;
	assert RAM(23090) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23090))))  severity failure;
	assert RAM(23091) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(23091))))  severity failure;
	assert RAM(23092) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(23092))))  severity failure;
	assert RAM(23093) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(23093))))  severity failure;
	assert RAM(23094) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23094))))  severity failure;
	assert RAM(23095) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(23095))))  severity failure;
	assert RAM(23096) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23096))))  severity failure;
	assert RAM(23097) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23097))))  severity failure;
	assert RAM(23098) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23098))))  severity failure;
	assert RAM(23099) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23099))))  severity failure;
	assert RAM(23100) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23100))))  severity failure;
	assert RAM(23101) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(23101))))  severity failure;
	assert RAM(23102) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23102))))  severity failure;
	assert RAM(23103) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23103))))  severity failure;
	assert RAM(23104) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(23104))))  severity failure;
	assert RAM(23105) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23105))))  severity failure;
	assert RAM(23106) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23106))))  severity failure;
	assert RAM(23107) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23107))))  severity failure;
	assert RAM(23108) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23108))))  severity failure;
	assert RAM(23109) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23109))))  severity failure;
	assert RAM(23110) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23110))))  severity failure;
	assert RAM(23111) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23111))))  severity failure;
	assert RAM(23112) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(23112))))  severity failure;
	assert RAM(23113) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(23113))))  severity failure;
	assert RAM(23114) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(23114))))  severity failure;
	assert RAM(23115) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23115))))  severity failure;
	assert RAM(23116) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23116))))  severity failure;
	assert RAM(23117) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23117))))  severity failure;
	assert RAM(23118) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23118))))  severity failure;
	assert RAM(23119) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(23119))))  severity failure;
	assert RAM(23120) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23120))))  severity failure;
	assert RAM(23121) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(23121))))  severity failure;
	assert RAM(23122) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23122))))  severity failure;
	assert RAM(23123) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(23123))))  severity failure;
	assert RAM(23124) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23124))))  severity failure;
	assert RAM(23125) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(23125))))  severity failure;
	assert RAM(23126) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23126))))  severity failure;
	assert RAM(23127) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23127))))  severity failure;
	assert RAM(23128) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23128))))  severity failure;
	assert RAM(23129) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(23129))))  severity failure;
	assert RAM(23130) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23130))))  severity failure;
	assert RAM(23131) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23131))))  severity failure;
	assert RAM(23132) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23132))))  severity failure;
	assert RAM(23133) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23133))))  severity failure;
	assert RAM(23134) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(23134))))  severity failure;
	assert RAM(23135) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(23135))))  severity failure;
	assert RAM(23136) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(23136))))  severity failure;
	assert RAM(23137) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(23137))))  severity failure;
	assert RAM(23138) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(23138))))  severity failure;
	assert RAM(23139) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(23139))))  severity failure;
	assert RAM(23140) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(23140))))  severity failure;
	assert RAM(23141) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(23141))))  severity failure;
	assert RAM(23142) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23142))))  severity failure;
	assert RAM(23143) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(23143))))  severity failure;
	assert RAM(23144) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23144))))  severity failure;
	assert RAM(23145) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(23145))))  severity failure;
	assert RAM(23146) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(23146))))  severity failure;
	assert RAM(23147) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23147))))  severity failure;
	assert RAM(23148) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23148))))  severity failure;
	assert RAM(23149) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(23149))))  severity failure;
	assert RAM(23150) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23150))))  severity failure;
	assert RAM(23151) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23151))))  severity failure;
	assert RAM(23152) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(23152))))  severity failure;
	assert RAM(23153) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23153))))  severity failure;
	assert RAM(23154) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23154))))  severity failure;
	assert RAM(23155) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(23155))))  severity failure;
	assert RAM(23156) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23156))))  severity failure;
	assert RAM(23157) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23157))))  severity failure;
	assert RAM(23158) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23158))))  severity failure;
	assert RAM(23159) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(23159))))  severity failure;
	assert RAM(23160) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23160))))  severity failure;
	assert RAM(23161) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23161))))  severity failure;
	assert RAM(23162) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23162))))  severity failure;
	assert RAM(23163) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23163))))  severity failure;
	assert RAM(23164) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(23164))))  severity failure;
	assert RAM(23165) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23165))))  severity failure;
	assert RAM(23166) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(23166))))  severity failure;
	assert RAM(23167) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23167))))  severity failure;
	assert RAM(23168) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(23168))))  severity failure;
	assert RAM(23169) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23169))))  severity failure;
	assert RAM(23170) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23170))))  severity failure;
	assert RAM(23171) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23171))))  severity failure;
	assert RAM(23172) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23172))))  severity failure;
	assert RAM(23173) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(23173))))  severity failure;
	assert RAM(23174) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23174))))  severity failure;
	assert RAM(23175) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(23175))))  severity failure;
	assert RAM(23176) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(23176))))  severity failure;
	assert RAM(23177) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23177))))  severity failure;
	assert RAM(23178) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23178))))  severity failure;
	assert RAM(23179) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23179))))  severity failure;
	assert RAM(23180) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23180))))  severity failure;
	assert RAM(23181) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(23181))))  severity failure;
	assert RAM(23182) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23182))))  severity failure;
	assert RAM(23183) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23183))))  severity failure;
	assert RAM(23184) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23184))))  severity failure;
	assert RAM(23185) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23185))))  severity failure;
	assert RAM(23186) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(23186))))  severity failure;
	assert RAM(23187) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23187))))  severity failure;
	assert RAM(23188) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(23188))))  severity failure;
	assert RAM(23189) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(23189))))  severity failure;
	assert RAM(23190) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(23190))))  severity failure;
	assert RAM(23191) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(23191))))  severity failure;
	assert RAM(23192) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(23192))))  severity failure;
	assert RAM(23193) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23193))))  severity failure;
	assert RAM(23194) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23194))))  severity failure;
	assert RAM(23195) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23195))))  severity failure;
	assert RAM(23196) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23196))))  severity failure;
	assert RAM(23197) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23197))))  severity failure;
	assert RAM(23198) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(23198))))  severity failure;
	assert RAM(23199) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(23199))))  severity failure;
	assert RAM(23200) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23200))))  severity failure;
	assert RAM(23201) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(23201))))  severity failure;
	assert RAM(23202) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23202))))  severity failure;
	assert RAM(23203) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(23203))))  severity failure;
	assert RAM(23204) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23204))))  severity failure;
	assert RAM(23205) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23205))))  severity failure;
	assert RAM(23206) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23206))))  severity failure;
	assert RAM(23207) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(23207))))  severity failure;
	assert RAM(23208) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(23208))))  severity failure;
	assert RAM(23209) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(23209))))  severity failure;
	assert RAM(23210) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23210))))  severity failure;
	assert RAM(23211) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(23211))))  severity failure;
	assert RAM(23212) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(23212))))  severity failure;
	assert RAM(23213) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23213))))  severity failure;
	assert RAM(23214) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23214))))  severity failure;
	assert RAM(23215) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23215))))  severity failure;
	assert RAM(23216) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23216))))  severity failure;
	assert RAM(23217) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(23217))))  severity failure;
	assert RAM(23218) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23218))))  severity failure;
	assert RAM(23219) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(23219))))  severity failure;
	assert RAM(23220) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(23220))))  severity failure;
	assert RAM(23221) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23221))))  severity failure;
	assert RAM(23222) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(23222))))  severity failure;
	assert RAM(23223) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(23223))))  severity failure;
	assert RAM(23224) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(23224))))  severity failure;
	assert RAM(23225) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23225))))  severity failure;
	assert RAM(23226) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(23226))))  severity failure;
	assert RAM(23227) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23227))))  severity failure;
	assert RAM(23228) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(23228))))  severity failure;
	assert RAM(23229) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(23229))))  severity failure;
	assert RAM(23230) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23230))))  severity failure;
	assert RAM(23231) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(23231))))  severity failure;
	assert RAM(23232) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(23232))))  severity failure;
	assert RAM(23233) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23233))))  severity failure;
	assert RAM(23234) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(23234))))  severity failure;
	assert RAM(23235) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23235))))  severity failure;
	assert RAM(23236) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(23236))))  severity failure;
	assert RAM(23237) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(23237))))  severity failure;
	assert RAM(23238) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23238))))  severity failure;
	assert RAM(23239) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(23239))))  severity failure;
	assert RAM(23240) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23240))))  severity failure;
	assert RAM(23241) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23241))))  severity failure;
	assert RAM(23242) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23242))))  severity failure;
	assert RAM(23243) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(23243))))  severity failure;
	assert RAM(23244) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23244))))  severity failure;
	assert RAM(23245) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(23245))))  severity failure;
	assert RAM(23246) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23246))))  severity failure;
	assert RAM(23247) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(23247))))  severity failure;
	assert RAM(23248) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23248))))  severity failure;
	assert RAM(23249) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23249))))  severity failure;
	assert RAM(23250) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23250))))  severity failure;
	assert RAM(23251) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23251))))  severity failure;
	assert RAM(23252) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23252))))  severity failure;
	assert RAM(23253) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(23253))))  severity failure;
	assert RAM(23254) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(23254))))  severity failure;
	assert RAM(23255) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23255))))  severity failure;
	assert RAM(23256) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(23256))))  severity failure;
	assert RAM(23257) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(23257))))  severity failure;
	assert RAM(23258) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(23258))))  severity failure;
	assert RAM(23259) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(23259))))  severity failure;
	assert RAM(23260) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23260))))  severity failure;
	assert RAM(23261) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23261))))  severity failure;
	assert RAM(23262) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23262))))  severity failure;
	assert RAM(23263) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23263))))  severity failure;
	assert RAM(23264) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23264))))  severity failure;
	assert RAM(23265) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(23265))))  severity failure;
	assert RAM(23266) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23266))))  severity failure;
	assert RAM(23267) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(23267))))  severity failure;
	assert RAM(23268) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23268))))  severity failure;
	assert RAM(23269) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23269))))  severity failure;
	assert RAM(23270) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23270))))  severity failure;
	assert RAM(23271) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23271))))  severity failure;
	assert RAM(23272) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(23272))))  severity failure;
	assert RAM(23273) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23273))))  severity failure;
	assert RAM(23274) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(23274))))  severity failure;
	assert RAM(23275) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23275))))  severity failure;
	assert RAM(23276) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(23276))))  severity failure;
	assert RAM(23277) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23277))))  severity failure;
	assert RAM(23278) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23278))))  severity failure;
	assert RAM(23279) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(23279))))  severity failure;
	assert RAM(23280) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23280))))  severity failure;
	assert RAM(23281) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(23281))))  severity failure;
	assert RAM(23282) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(23282))))  severity failure;
	assert RAM(23283) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23283))))  severity failure;
	assert RAM(23284) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23284))))  severity failure;
	assert RAM(23285) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23285))))  severity failure;
	assert RAM(23286) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(23286))))  severity failure;
	assert RAM(23287) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23287))))  severity failure;
	assert RAM(23288) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23288))))  severity failure;
	assert RAM(23289) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(23289))))  severity failure;
	assert RAM(23290) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23290))))  severity failure;
	assert RAM(23291) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(23291))))  severity failure;
	assert RAM(23292) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23292))))  severity failure;
	assert RAM(23293) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23293))))  severity failure;
	assert RAM(23294) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(23294))))  severity failure;
	assert RAM(23295) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23295))))  severity failure;
	assert RAM(23296) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23296))))  severity failure;
	assert RAM(23297) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(23297))))  severity failure;
	assert RAM(23298) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(23298))))  severity failure;
	assert RAM(23299) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23299))))  severity failure;
	assert RAM(23300) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(23300))))  severity failure;
	assert RAM(23301) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23301))))  severity failure;
	assert RAM(23302) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(23302))))  severity failure;
	assert RAM(23303) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(23303))))  severity failure;
	assert RAM(23304) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23304))))  severity failure;
	assert RAM(23305) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(23305))))  severity failure;
	assert RAM(23306) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(23306))))  severity failure;
	assert RAM(23307) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(23307))))  severity failure;
	assert RAM(23308) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23308))))  severity failure;
	assert RAM(23309) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(23309))))  severity failure;
	assert RAM(23310) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(23310))))  severity failure;
	assert RAM(23311) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(23311))))  severity failure;
	assert RAM(23312) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23312))))  severity failure;
	assert RAM(23313) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(23313))))  severity failure;
	assert RAM(23314) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23314))))  severity failure;
	assert RAM(23315) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23315))))  severity failure;
	assert RAM(23316) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23316))))  severity failure;
	assert RAM(23317) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23317))))  severity failure;
	assert RAM(23318) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23318))))  severity failure;
	assert RAM(23319) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23319))))  severity failure;
	assert RAM(23320) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(23320))))  severity failure;
	assert RAM(23321) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(23321))))  severity failure;
	assert RAM(23322) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(23322))))  severity failure;
	assert RAM(23323) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(23323))))  severity failure;
	assert RAM(23324) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23324))))  severity failure;
	assert RAM(23325) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23325))))  severity failure;
	assert RAM(23326) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(23326))))  severity failure;
	assert RAM(23327) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23327))))  severity failure;
	assert RAM(23328) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(23328))))  severity failure;
	assert RAM(23329) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(23329))))  severity failure;
	assert RAM(23330) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(23330))))  severity failure;
	assert RAM(23331) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23331))))  severity failure;
	assert RAM(23332) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23332))))  severity failure;
	assert RAM(23333) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23333))))  severity failure;
	assert RAM(23334) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23334))))  severity failure;
	assert RAM(23335) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23335))))  severity failure;
	assert RAM(23336) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(23336))))  severity failure;
	assert RAM(23337) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(23337))))  severity failure;
	assert RAM(23338) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(23338))))  severity failure;
	assert RAM(23339) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23339))))  severity failure;
	assert RAM(23340) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23340))))  severity failure;
	assert RAM(23341) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23341))))  severity failure;
	assert RAM(23342) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23342))))  severity failure;
	assert RAM(23343) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23343))))  severity failure;
	assert RAM(23344) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23344))))  severity failure;
	assert RAM(23345) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23345))))  severity failure;
	assert RAM(23346) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(23346))))  severity failure;
	assert RAM(23347) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(23347))))  severity failure;
	assert RAM(23348) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23348))))  severity failure;
	assert RAM(23349) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(23349))))  severity failure;
	assert RAM(23350) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23350))))  severity failure;
	assert RAM(23351) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23351))))  severity failure;
	assert RAM(23352) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(23352))))  severity failure;
	assert RAM(23353) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(23353))))  severity failure;
	assert RAM(23354) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23354))))  severity failure;
	assert RAM(23355) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(23355))))  severity failure;
	assert RAM(23356) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23356))))  severity failure;
	assert RAM(23357) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23357))))  severity failure;
	assert RAM(23358) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23358))))  severity failure;
	assert RAM(23359) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23359))))  severity failure;
	assert RAM(23360) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(23360))))  severity failure;
	assert RAM(23361) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(23361))))  severity failure;
	assert RAM(23362) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23362))))  severity failure;
	assert RAM(23363) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23363))))  severity failure;
	assert RAM(23364) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(23364))))  severity failure;
	assert RAM(23365) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(23365))))  severity failure;
	assert RAM(23366) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23366))))  severity failure;
	assert RAM(23367) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23367))))  severity failure;
	assert RAM(23368) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23368))))  severity failure;
	assert RAM(23369) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(23369))))  severity failure;
	assert RAM(23370) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(23370))))  severity failure;
	assert RAM(23371) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(23371))))  severity failure;
	assert RAM(23372) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23372))))  severity failure;
	assert RAM(23373) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(23373))))  severity failure;
	assert RAM(23374) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(23374))))  severity failure;
	assert RAM(23375) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(23375))))  severity failure;
	assert RAM(23376) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23376))))  severity failure;
	assert RAM(23377) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23377))))  severity failure;
	assert RAM(23378) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(23378))))  severity failure;
	assert RAM(23379) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(23379))))  severity failure;
	assert RAM(23380) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(23380))))  severity failure;
	assert RAM(23381) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23381))))  severity failure;
	assert RAM(23382) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23382))))  severity failure;
	assert RAM(23383) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(23383))))  severity failure;
	assert RAM(23384) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23384))))  severity failure;
	assert RAM(23385) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23385))))  severity failure;
	assert RAM(23386) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(23386))))  severity failure;
	assert RAM(23387) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23387))))  severity failure;
	assert RAM(23388) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23388))))  severity failure;
	assert RAM(23389) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(23389))))  severity failure;
	assert RAM(23390) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(23390))))  severity failure;
	assert RAM(23391) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(23391))))  severity failure;
	assert RAM(23392) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23392))))  severity failure;
	assert RAM(23393) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23393))))  severity failure;
	assert RAM(23394) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23394))))  severity failure;
	assert RAM(23395) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23395))))  severity failure;
	assert RAM(23396) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23396))))  severity failure;
	assert RAM(23397) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23397))))  severity failure;
	assert RAM(23398) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(23398))))  severity failure;
	assert RAM(23399) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23399))))  severity failure;
	assert RAM(23400) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(23400))))  severity failure;
	assert RAM(23401) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23401))))  severity failure;
	assert RAM(23402) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23402))))  severity failure;
	assert RAM(23403) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(23403))))  severity failure;
	assert RAM(23404) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23404))))  severity failure;
	assert RAM(23405) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(23405))))  severity failure;
	assert RAM(23406) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23406))))  severity failure;
	assert RAM(23407) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23407))))  severity failure;
	assert RAM(23408) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(23408))))  severity failure;
	assert RAM(23409) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23409))))  severity failure;
	assert RAM(23410) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23410))))  severity failure;
	assert RAM(23411) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23411))))  severity failure;
	assert RAM(23412) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23412))))  severity failure;
	assert RAM(23413) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(23413))))  severity failure;
	assert RAM(23414) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23414))))  severity failure;
	assert RAM(23415) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23415))))  severity failure;
	assert RAM(23416) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(23416))))  severity failure;
	assert RAM(23417) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23417))))  severity failure;
	assert RAM(23418) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(23418))))  severity failure;
	assert RAM(23419) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(23419))))  severity failure;
	assert RAM(23420) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(23420))))  severity failure;
	assert RAM(23421) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(23421))))  severity failure;
	assert RAM(23422) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(23422))))  severity failure;
	assert RAM(23423) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23423))))  severity failure;
	assert RAM(23424) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23424))))  severity failure;
	assert RAM(23425) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(23425))))  severity failure;
	assert RAM(23426) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(23426))))  severity failure;
	assert RAM(23427) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(23427))))  severity failure;
	assert RAM(23428) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23428))))  severity failure;
	assert RAM(23429) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(23429))))  severity failure;
	assert RAM(23430) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23430))))  severity failure;
	assert RAM(23431) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23431))))  severity failure;
	assert RAM(23432) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(23432))))  severity failure;
	assert RAM(23433) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23433))))  severity failure;
	assert RAM(23434) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(23434))))  severity failure;
	assert RAM(23435) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(23435))))  severity failure;
	assert RAM(23436) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(23436))))  severity failure;
	assert RAM(23437) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23437))))  severity failure;
	assert RAM(23438) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23438))))  severity failure;
	assert RAM(23439) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(23439))))  severity failure;
	assert RAM(23440) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23440))))  severity failure;
	assert RAM(23441) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23441))))  severity failure;
	assert RAM(23442) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(23442))))  severity failure;
	assert RAM(23443) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(23443))))  severity failure;
	assert RAM(23444) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23444))))  severity failure;
	assert RAM(23445) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23445))))  severity failure;
	assert RAM(23446) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23446))))  severity failure;
	assert RAM(23447) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(23447))))  severity failure;
	assert RAM(23448) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(23448))))  severity failure;
	assert RAM(23449) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(23449))))  severity failure;
	assert RAM(23450) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23450))))  severity failure;
	assert RAM(23451) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23451))))  severity failure;
	assert RAM(23452) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(23452))))  severity failure;
	assert RAM(23453) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23453))))  severity failure;
	assert RAM(23454) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23454))))  severity failure;
	assert RAM(23455) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23455))))  severity failure;
	assert RAM(23456) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(23456))))  severity failure;
	assert RAM(23457) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(23457))))  severity failure;
	assert RAM(23458) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(23458))))  severity failure;
	assert RAM(23459) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(23459))))  severity failure;
	assert RAM(23460) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23460))))  severity failure;
	assert RAM(23461) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23461))))  severity failure;
	assert RAM(23462) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(23462))))  severity failure;
	assert RAM(23463) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(23463))))  severity failure;
	assert RAM(23464) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23464))))  severity failure;
	assert RAM(23465) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(23465))))  severity failure;
	assert RAM(23466) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23466))))  severity failure;
	assert RAM(23467) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23467))))  severity failure;
	assert RAM(23468) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(23468))))  severity failure;
	assert RAM(23469) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(23469))))  severity failure;
	assert RAM(23470) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(23470))))  severity failure;
	assert RAM(23471) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23471))))  severity failure;
	assert RAM(23472) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23472))))  severity failure;
	assert RAM(23473) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(23473))))  severity failure;
	assert RAM(23474) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(23474))))  severity failure;
	assert RAM(23475) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(23475))))  severity failure;
	assert RAM(23476) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(23476))))  severity failure;
	assert RAM(23477) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23477))))  severity failure;
	assert RAM(23478) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(23478))))  severity failure;
	assert RAM(23479) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(23479))))  severity failure;
	assert RAM(23480) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(23480))))  severity failure;
	assert RAM(23481) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23481))))  severity failure;
	assert RAM(23482) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(23482))))  severity failure;
	assert RAM(23483) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(23483))))  severity failure;
	assert RAM(23484) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(23484))))  severity failure;
	assert RAM(23485) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(23485))))  severity failure;
	assert RAM(23486) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(23486))))  severity failure;
	assert RAM(23487) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(23487))))  severity failure;
	assert RAM(23488) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23488))))  severity failure;
	assert RAM(23489) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23489))))  severity failure;
	assert RAM(23490) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23490))))  severity failure;
	assert RAM(23491) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23491))))  severity failure;
	assert RAM(23492) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23492))))  severity failure;
	assert RAM(23493) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(23493))))  severity failure;
	assert RAM(23494) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23494))))  severity failure;
	assert RAM(23495) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(23495))))  severity failure;
	assert RAM(23496) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(23496))))  severity failure;
	assert RAM(23497) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23497))))  severity failure;
	assert RAM(23498) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23498))))  severity failure;
	assert RAM(23499) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(23499))))  severity failure;
	assert RAM(23500) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23500))))  severity failure;
	assert RAM(23501) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23501))))  severity failure;
	assert RAM(23502) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(23502))))  severity failure;
	assert RAM(23503) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23503))))  severity failure;
	assert RAM(23504) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23504))))  severity failure;
	assert RAM(23505) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23505))))  severity failure;
	assert RAM(23506) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23506))))  severity failure;
	assert RAM(23507) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(23507))))  severity failure;
	assert RAM(23508) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(23508))))  severity failure;
	assert RAM(23509) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(23509))))  severity failure;
	assert RAM(23510) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23510))))  severity failure;
	assert RAM(23511) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23511))))  severity failure;
	assert RAM(23512) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(23512))))  severity failure;
	assert RAM(23513) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23513))))  severity failure;
	assert RAM(23514) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(23514))))  severity failure;
	assert RAM(23515) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(23515))))  severity failure;
	assert RAM(23516) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23516))))  severity failure;
	assert RAM(23517) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(23517))))  severity failure;
	assert RAM(23518) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23518))))  severity failure;
	assert RAM(23519) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23519))))  severity failure;
	assert RAM(23520) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(23520))))  severity failure;
	assert RAM(23521) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(23521))))  severity failure;
	assert RAM(23522) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(23522))))  severity failure;
	assert RAM(23523) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23523))))  severity failure;
	assert RAM(23524) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(23524))))  severity failure;
	assert RAM(23525) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(23525))))  severity failure;
	assert RAM(23526) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(23526))))  severity failure;
	assert RAM(23527) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23527))))  severity failure;
	assert RAM(23528) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(23528))))  severity failure;
	assert RAM(23529) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23529))))  severity failure;
	assert RAM(23530) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23530))))  severity failure;
	assert RAM(23531) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(23531))))  severity failure;
	assert RAM(23532) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23532))))  severity failure;
	assert RAM(23533) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23533))))  severity failure;
	assert RAM(23534) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(23534))))  severity failure;
	assert RAM(23535) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(23535))))  severity failure;
	assert RAM(23536) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23536))))  severity failure;
	assert RAM(23537) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23537))))  severity failure;
	assert RAM(23538) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23538))))  severity failure;
	assert RAM(23539) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(23539))))  severity failure;
	assert RAM(23540) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(23540))))  severity failure;
	assert RAM(23541) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(23541))))  severity failure;
	assert RAM(23542) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23542))))  severity failure;
	assert RAM(23543) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23543))))  severity failure;
	assert RAM(23544) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23544))))  severity failure;
	assert RAM(23545) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23545))))  severity failure;
	assert RAM(23546) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23546))))  severity failure;
	assert RAM(23547) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(23547))))  severity failure;
	assert RAM(23548) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23548))))  severity failure;
	assert RAM(23549) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(23549))))  severity failure;
	assert RAM(23550) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23550))))  severity failure;
	assert RAM(23551) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23551))))  severity failure;
	assert RAM(23552) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23552))))  severity failure;
	assert RAM(23553) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23553))))  severity failure;
	assert RAM(23554) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23554))))  severity failure;
	assert RAM(23555) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23555))))  severity failure;
	assert RAM(23556) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23556))))  severity failure;
	assert RAM(23557) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(23557))))  severity failure;
	assert RAM(23558) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(23558))))  severity failure;
	assert RAM(23559) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23559))))  severity failure;
	assert RAM(23560) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(23560))))  severity failure;
	assert RAM(23561) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23561))))  severity failure;
	assert RAM(23562) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23562))))  severity failure;
	assert RAM(23563) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23563))))  severity failure;
	assert RAM(23564) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23564))))  severity failure;
	assert RAM(23565) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23565))))  severity failure;
	assert RAM(23566) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23566))))  severity failure;
	assert RAM(23567) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(23567))))  severity failure;
	assert RAM(23568) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(23568))))  severity failure;
	assert RAM(23569) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23569))))  severity failure;
	assert RAM(23570) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23570))))  severity failure;
	assert RAM(23571) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23571))))  severity failure;
	assert RAM(23572) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23572))))  severity failure;
	assert RAM(23573) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(23573))))  severity failure;
	assert RAM(23574) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23574))))  severity failure;
	assert RAM(23575) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23575))))  severity failure;
	assert RAM(23576) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23576))))  severity failure;
	assert RAM(23577) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(23577))))  severity failure;
	assert RAM(23578) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23578))))  severity failure;
	assert RAM(23579) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(23579))))  severity failure;
	assert RAM(23580) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(23580))))  severity failure;
	assert RAM(23581) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23581))))  severity failure;
	assert RAM(23582) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23582))))  severity failure;
	assert RAM(23583) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23583))))  severity failure;
	assert RAM(23584) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(23584))))  severity failure;
	assert RAM(23585) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23585))))  severity failure;
	assert RAM(23586) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23586))))  severity failure;
	assert RAM(23587) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23587))))  severity failure;
	assert RAM(23588) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23588))))  severity failure;
	assert RAM(23589) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23589))))  severity failure;
	assert RAM(23590) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(23590))))  severity failure;
	assert RAM(23591) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23591))))  severity failure;
	assert RAM(23592) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23592))))  severity failure;
	assert RAM(23593) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(23593))))  severity failure;
	assert RAM(23594) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(23594))))  severity failure;
	assert RAM(23595) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(23595))))  severity failure;
	assert RAM(23596) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23596))))  severity failure;
	assert RAM(23597) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(23597))))  severity failure;
	assert RAM(23598) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23598))))  severity failure;
	assert RAM(23599) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(23599))))  severity failure;
	assert RAM(23600) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23600))))  severity failure;
	assert RAM(23601) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(23601))))  severity failure;
	assert RAM(23602) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23602))))  severity failure;
	assert RAM(23603) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23603))))  severity failure;
	assert RAM(23604) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23604))))  severity failure;
	assert RAM(23605) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(23605))))  severity failure;
	assert RAM(23606) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23606))))  severity failure;
	assert RAM(23607) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23607))))  severity failure;
	assert RAM(23608) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23608))))  severity failure;
	assert RAM(23609) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23609))))  severity failure;
	assert RAM(23610) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(23610))))  severity failure;
	assert RAM(23611) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(23611))))  severity failure;
	assert RAM(23612) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23612))))  severity failure;
	assert RAM(23613) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(23613))))  severity failure;
	assert RAM(23614) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23614))))  severity failure;
	assert RAM(23615) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23615))))  severity failure;
	assert RAM(23616) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23616))))  severity failure;
	assert RAM(23617) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(23617))))  severity failure;
	assert RAM(23618) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(23618))))  severity failure;
	assert RAM(23619) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23619))))  severity failure;
	assert RAM(23620) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23620))))  severity failure;
	assert RAM(23621) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23621))))  severity failure;
	assert RAM(23622) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(23622))))  severity failure;
	assert RAM(23623) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(23623))))  severity failure;
	assert RAM(23624) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23624))))  severity failure;
	assert RAM(23625) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23625))))  severity failure;
	assert RAM(23626) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23626))))  severity failure;
	assert RAM(23627) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23627))))  severity failure;
	assert RAM(23628) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23628))))  severity failure;
	assert RAM(23629) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(23629))))  severity failure;
	assert RAM(23630) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23630))))  severity failure;
	assert RAM(23631) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23631))))  severity failure;
	assert RAM(23632) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(23632))))  severity failure;
	assert RAM(23633) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23633))))  severity failure;
	assert RAM(23634) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23634))))  severity failure;
	assert RAM(23635) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23635))))  severity failure;
	assert RAM(23636) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(23636))))  severity failure;
	assert RAM(23637) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23637))))  severity failure;
	assert RAM(23638) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(23638))))  severity failure;
	assert RAM(23639) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(23639))))  severity failure;
	assert RAM(23640) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23640))))  severity failure;
	assert RAM(23641) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23641))))  severity failure;
	assert RAM(23642) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23642))))  severity failure;
	assert RAM(23643) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(23643))))  severity failure;
	assert RAM(23644) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(23644))))  severity failure;
	assert RAM(23645) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(23645))))  severity failure;
	assert RAM(23646) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23646))))  severity failure;
	assert RAM(23647) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(23647))))  severity failure;
	assert RAM(23648) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(23648))))  severity failure;
	assert RAM(23649) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(23649))))  severity failure;
	assert RAM(23650) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23650))))  severity failure;
	assert RAM(23651) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23651))))  severity failure;
	assert RAM(23652) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(23652))))  severity failure;
	assert RAM(23653) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23653))))  severity failure;
	assert RAM(23654) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23654))))  severity failure;
	assert RAM(23655) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23655))))  severity failure;
	assert RAM(23656) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(23656))))  severity failure;
	assert RAM(23657) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23657))))  severity failure;
	assert RAM(23658) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23658))))  severity failure;
	assert RAM(23659) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(23659))))  severity failure;
	assert RAM(23660) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(23660))))  severity failure;
	assert RAM(23661) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(23661))))  severity failure;
	assert RAM(23662) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23662))))  severity failure;
	assert RAM(23663) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(23663))))  severity failure;
	assert RAM(23664) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(23664))))  severity failure;
	assert RAM(23665) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23665))))  severity failure;
	assert RAM(23666) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(23666))))  severity failure;
	assert RAM(23667) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(23667))))  severity failure;
	assert RAM(23668) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23668))))  severity failure;
	assert RAM(23669) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(23669))))  severity failure;
	assert RAM(23670) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23670))))  severity failure;
	assert RAM(23671) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23671))))  severity failure;
	assert RAM(23672) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23672))))  severity failure;
	assert RAM(23673) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(23673))))  severity failure;
	assert RAM(23674) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(23674))))  severity failure;
	assert RAM(23675) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23675))))  severity failure;
	assert RAM(23676) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(23676))))  severity failure;
	assert RAM(23677) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(23677))))  severity failure;
	assert RAM(23678) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23678))))  severity failure;
	assert RAM(23679) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23679))))  severity failure;
	assert RAM(23680) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(23680))))  severity failure;
	assert RAM(23681) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(23681))))  severity failure;
	assert RAM(23682) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(23682))))  severity failure;
	assert RAM(23683) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23683))))  severity failure;
	assert RAM(23684) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(23684))))  severity failure;
	assert RAM(23685) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23685))))  severity failure;
	assert RAM(23686) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23686))))  severity failure;
	assert RAM(23687) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(23687))))  severity failure;
	assert RAM(23688) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23688))))  severity failure;
	assert RAM(23689) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(23689))))  severity failure;
	assert RAM(23690) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23690))))  severity failure;
	assert RAM(23691) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23691))))  severity failure;
	assert RAM(23692) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(23692))))  severity failure;
	assert RAM(23693) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(23693))))  severity failure;
	assert RAM(23694) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(23694))))  severity failure;
	assert RAM(23695) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23695))))  severity failure;
	assert RAM(23696) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(23696))))  severity failure;
	assert RAM(23697) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(23697))))  severity failure;
	assert RAM(23698) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23698))))  severity failure;
	assert RAM(23699) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(23699))))  severity failure;
	assert RAM(23700) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(23700))))  severity failure;
	assert RAM(23701) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(23701))))  severity failure;
	assert RAM(23702) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23702))))  severity failure;
	assert RAM(23703) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23703))))  severity failure;
	assert RAM(23704) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(23704))))  severity failure;
	assert RAM(23705) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23705))))  severity failure;
	assert RAM(23706) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(23706))))  severity failure;
	assert RAM(23707) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(23707))))  severity failure;
	assert RAM(23708) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(23708))))  severity failure;
	assert RAM(23709) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23709))))  severity failure;
	assert RAM(23710) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(23710))))  severity failure;
	assert RAM(23711) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(23711))))  severity failure;
	assert RAM(23712) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23712))))  severity failure;
	assert RAM(23713) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(23713))))  severity failure;
	assert RAM(23714) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23714))))  severity failure;
	assert RAM(23715) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(23715))))  severity failure;
	assert RAM(23716) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(23716))))  severity failure;
	assert RAM(23717) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(23717))))  severity failure;
	assert RAM(23718) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23718))))  severity failure;
	assert RAM(23719) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(23719))))  severity failure;
	assert RAM(23720) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(23720))))  severity failure;
	assert RAM(23721) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23721))))  severity failure;
	assert RAM(23722) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23722))))  severity failure;
	assert RAM(23723) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23723))))  severity failure;
	assert RAM(23724) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23724))))  severity failure;
	assert RAM(23725) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23725))))  severity failure;
	assert RAM(23726) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23726))))  severity failure;
	assert RAM(23727) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23727))))  severity failure;
	assert RAM(23728) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23728))))  severity failure;
	assert RAM(23729) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23729))))  severity failure;
	assert RAM(23730) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(23730))))  severity failure;
	assert RAM(23731) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23731))))  severity failure;
	assert RAM(23732) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(23732))))  severity failure;
	assert RAM(23733) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23733))))  severity failure;
	assert RAM(23734) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23734))))  severity failure;
	assert RAM(23735) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(23735))))  severity failure;
	assert RAM(23736) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(23736))))  severity failure;
	assert RAM(23737) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23737))))  severity failure;
	assert RAM(23738) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(23738))))  severity failure;
	assert RAM(23739) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(23739))))  severity failure;
	assert RAM(23740) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23740))))  severity failure;
	assert RAM(23741) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23741))))  severity failure;
	assert RAM(23742) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(23742))))  severity failure;
	assert RAM(23743) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23743))))  severity failure;
	assert RAM(23744) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(23744))))  severity failure;
	assert RAM(23745) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23745))))  severity failure;
	assert RAM(23746) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23746))))  severity failure;
	assert RAM(23747) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(23747))))  severity failure;
	assert RAM(23748) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23748))))  severity failure;
	assert RAM(23749) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(23749))))  severity failure;
	assert RAM(23750) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23750))))  severity failure;
	assert RAM(23751) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23751))))  severity failure;
	assert RAM(23752) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23752))))  severity failure;
	assert RAM(23753) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(23753))))  severity failure;
	assert RAM(23754) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23754))))  severity failure;
	assert RAM(23755) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(23755))))  severity failure;
	assert RAM(23756) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23756))))  severity failure;
	assert RAM(23757) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23757))))  severity failure;
	assert RAM(23758) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23758))))  severity failure;
	assert RAM(23759) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(23759))))  severity failure;
	assert RAM(23760) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23760))))  severity failure;
	assert RAM(23761) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23761))))  severity failure;
	assert RAM(23762) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23762))))  severity failure;
	assert RAM(23763) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23763))))  severity failure;
	assert RAM(23764) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23764))))  severity failure;
	assert RAM(23765) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23765))))  severity failure;
	assert RAM(23766) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(23766))))  severity failure;
	assert RAM(23767) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23767))))  severity failure;
	assert RAM(23768) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23768))))  severity failure;
	assert RAM(23769) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23769))))  severity failure;
	assert RAM(23770) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(23770))))  severity failure;
	assert RAM(23771) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(23771))))  severity failure;
	assert RAM(23772) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23772))))  severity failure;
	assert RAM(23773) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23773))))  severity failure;
	assert RAM(23774) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23774))))  severity failure;
	assert RAM(23775) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23775))))  severity failure;
	assert RAM(23776) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(23776))))  severity failure;
	assert RAM(23777) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(23777))))  severity failure;
	assert RAM(23778) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(23778))))  severity failure;
	assert RAM(23779) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(23779))))  severity failure;
	assert RAM(23780) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(23780))))  severity failure;
	assert RAM(23781) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(23781))))  severity failure;
	assert RAM(23782) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(23782))))  severity failure;
	assert RAM(23783) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23783))))  severity failure;
	assert RAM(23784) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(23784))))  severity failure;
	assert RAM(23785) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(23785))))  severity failure;
	assert RAM(23786) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23786))))  severity failure;
	assert RAM(23787) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23787))))  severity failure;
	assert RAM(23788) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23788))))  severity failure;
	assert RAM(23789) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(23789))))  severity failure;
	assert RAM(23790) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23790))))  severity failure;
	assert RAM(23791) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23791))))  severity failure;
	assert RAM(23792) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23792))))  severity failure;
	assert RAM(23793) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(23793))))  severity failure;
	assert RAM(23794) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(23794))))  severity failure;
	assert RAM(23795) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(23795))))  severity failure;
	assert RAM(23796) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23796))))  severity failure;
	assert RAM(23797) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23797))))  severity failure;
	assert RAM(23798) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23798))))  severity failure;
	assert RAM(23799) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23799))))  severity failure;
	assert RAM(23800) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(23800))))  severity failure;
	assert RAM(23801) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(23801))))  severity failure;
	assert RAM(23802) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(23802))))  severity failure;
	assert RAM(23803) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23803))))  severity failure;
	assert RAM(23804) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23804))))  severity failure;
	assert RAM(23805) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23805))))  severity failure;
	assert RAM(23806) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23806))))  severity failure;
	assert RAM(23807) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23807))))  severity failure;
	assert RAM(23808) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(23808))))  severity failure;
	assert RAM(23809) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(23809))))  severity failure;
	assert RAM(23810) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23810))))  severity failure;
	assert RAM(23811) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23811))))  severity failure;
	assert RAM(23812) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23812))))  severity failure;
	assert RAM(23813) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23813))))  severity failure;
	assert RAM(23814) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23814))))  severity failure;
	assert RAM(23815) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(23815))))  severity failure;
	assert RAM(23816) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23816))))  severity failure;
	assert RAM(23817) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23817))))  severity failure;
	assert RAM(23818) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23818))))  severity failure;
	assert RAM(23819) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(23819))))  severity failure;
	assert RAM(23820) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23820))))  severity failure;
	assert RAM(23821) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23821))))  severity failure;
	assert RAM(23822) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(23822))))  severity failure;
	assert RAM(23823) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23823))))  severity failure;
	assert RAM(23824) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23824))))  severity failure;
	assert RAM(23825) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(23825))))  severity failure;
	assert RAM(23826) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23826))))  severity failure;
	assert RAM(23827) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(23827))))  severity failure;
	assert RAM(23828) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(23828))))  severity failure;
	assert RAM(23829) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23829))))  severity failure;
	assert RAM(23830) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23830))))  severity failure;
	assert RAM(23831) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(23831))))  severity failure;
	assert RAM(23832) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(23832))))  severity failure;
	assert RAM(23833) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23833))))  severity failure;
	assert RAM(23834) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23834))))  severity failure;
	assert RAM(23835) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23835))))  severity failure;
	assert RAM(23836) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(23836))))  severity failure;
	assert RAM(23837) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(23837))))  severity failure;
	assert RAM(23838) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(23838))))  severity failure;
	assert RAM(23839) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23839))))  severity failure;
	assert RAM(23840) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(23840))))  severity failure;
	assert RAM(23841) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(23841))))  severity failure;
	assert RAM(23842) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23842))))  severity failure;
	assert RAM(23843) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23843))))  severity failure;
	assert RAM(23844) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(23844))))  severity failure;
	assert RAM(23845) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(23845))))  severity failure;
	assert RAM(23846) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23846))))  severity failure;
	assert RAM(23847) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23847))))  severity failure;
	assert RAM(23848) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23848))))  severity failure;
	assert RAM(23849) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(23849))))  severity failure;
	assert RAM(23850) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23850))))  severity failure;
	assert RAM(23851) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(23851))))  severity failure;
	assert RAM(23852) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(23852))))  severity failure;
	assert RAM(23853) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(23853))))  severity failure;
	assert RAM(23854) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(23854))))  severity failure;
	assert RAM(23855) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23855))))  severity failure;
	assert RAM(23856) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23856))))  severity failure;
	assert RAM(23857) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(23857))))  severity failure;
	assert RAM(23858) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23858))))  severity failure;
	assert RAM(23859) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(23859))))  severity failure;
	assert RAM(23860) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(23860))))  severity failure;
	assert RAM(23861) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(23861))))  severity failure;
	assert RAM(23862) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(23862))))  severity failure;
	assert RAM(23863) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(23863))))  severity failure;
	assert RAM(23864) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23864))))  severity failure;
	assert RAM(23865) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23865))))  severity failure;
	assert RAM(23866) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23866))))  severity failure;
	assert RAM(23867) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(23867))))  severity failure;
	assert RAM(23868) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23868))))  severity failure;
	assert RAM(23869) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23869))))  severity failure;
	assert RAM(23870) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(23870))))  severity failure;
	assert RAM(23871) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23871))))  severity failure;
	assert RAM(23872) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(23872))))  severity failure;
	assert RAM(23873) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(23873))))  severity failure;
	assert RAM(23874) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(23874))))  severity failure;
	assert RAM(23875) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(23875))))  severity failure;
	assert RAM(23876) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(23876))))  severity failure;
	assert RAM(23877) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(23877))))  severity failure;
	assert RAM(23878) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(23878))))  severity failure;
	assert RAM(23879) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(23879))))  severity failure;
	assert RAM(23880) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23880))))  severity failure;
	assert RAM(23881) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23881))))  severity failure;
	assert RAM(23882) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23882))))  severity failure;
	assert RAM(23883) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(23883))))  severity failure;
	assert RAM(23884) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23884))))  severity failure;
	assert RAM(23885) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23885))))  severity failure;
	assert RAM(23886) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(23886))))  severity failure;
	assert RAM(23887) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23887))))  severity failure;
	assert RAM(23888) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23888))))  severity failure;
	assert RAM(23889) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23889))))  severity failure;
	assert RAM(23890) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(23890))))  severity failure;
	assert RAM(23891) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23891))))  severity failure;
	assert RAM(23892) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(23892))))  severity failure;
	assert RAM(23893) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23893))))  severity failure;
	assert RAM(23894) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(23894))))  severity failure;
	assert RAM(23895) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23895))))  severity failure;
	assert RAM(23896) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23896))))  severity failure;
	assert RAM(23897) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23897))))  severity failure;
	assert RAM(23898) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(23898))))  severity failure;
	assert RAM(23899) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23899))))  severity failure;
	assert RAM(23900) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23900))))  severity failure;
	assert RAM(23901) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23901))))  severity failure;
	assert RAM(23902) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(23902))))  severity failure;
	assert RAM(23903) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(23903))))  severity failure;
	assert RAM(23904) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(23904))))  severity failure;
	assert RAM(23905) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(23905))))  severity failure;
	assert RAM(23906) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23906))))  severity failure;
	assert RAM(23907) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(23907))))  severity failure;
	assert RAM(23908) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(23908))))  severity failure;
	assert RAM(23909) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23909))))  severity failure;
	assert RAM(23910) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23910))))  severity failure;
	assert RAM(23911) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23911))))  severity failure;
	assert RAM(23912) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(23912))))  severity failure;
	assert RAM(23913) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23913))))  severity failure;
	assert RAM(23914) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23914))))  severity failure;
	assert RAM(23915) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(23915))))  severity failure;
	assert RAM(23916) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23916))))  severity failure;
	assert RAM(23917) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23917))))  severity failure;
	assert RAM(23918) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(23918))))  severity failure;
	assert RAM(23919) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(23919))))  severity failure;
	assert RAM(23920) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(23920))))  severity failure;
	assert RAM(23921) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23921))))  severity failure;
	assert RAM(23922) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23922))))  severity failure;
	assert RAM(23923) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23923))))  severity failure;
	assert RAM(23924) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(23924))))  severity failure;
	assert RAM(23925) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(23925))))  severity failure;
	assert RAM(23926) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(23926))))  severity failure;
	assert RAM(23927) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23927))))  severity failure;
	assert RAM(23928) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23928))))  severity failure;
	assert RAM(23929) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(23929))))  severity failure;
	assert RAM(23930) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23930))))  severity failure;
	assert RAM(23931) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23931))))  severity failure;
	assert RAM(23932) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23932))))  severity failure;
	assert RAM(23933) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23933))))  severity failure;
	assert RAM(23934) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(23934))))  severity failure;
	assert RAM(23935) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23935))))  severity failure;
	assert RAM(23936) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23936))))  severity failure;
	assert RAM(23937) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23937))))  severity failure;
	assert RAM(23938) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(23938))))  severity failure;
	assert RAM(23939) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(23939))))  severity failure;
	assert RAM(23940) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23940))))  severity failure;
	assert RAM(23941) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(23941))))  severity failure;
	assert RAM(23942) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23942))))  severity failure;
	assert RAM(23943) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23943))))  severity failure;
	assert RAM(23944) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23944))))  severity failure;
	assert RAM(23945) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23945))))  severity failure;
	assert RAM(23946) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(23946))))  severity failure;
	assert RAM(23947) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(23947))))  severity failure;
	assert RAM(23948) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(23948))))  severity failure;
	assert RAM(23949) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23949))))  severity failure;
	assert RAM(23950) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(23950))))  severity failure;
	assert RAM(23951) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(23951))))  severity failure;
	assert RAM(23952) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23952))))  severity failure;
	assert RAM(23953) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(23953))))  severity failure;
	assert RAM(23954) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(23954))))  severity failure;
	assert RAM(23955) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(23955))))  severity failure;
	assert RAM(23956) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(23956))))  severity failure;
	assert RAM(23957) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23957))))  severity failure;
	assert RAM(23958) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23958))))  severity failure;
	assert RAM(23959) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(23959))))  severity failure;
	assert RAM(23960) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(23960))))  severity failure;
	assert RAM(23961) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23961))))  severity failure;
	assert RAM(23962) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(23962))))  severity failure;
	assert RAM(23963) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23963))))  severity failure;
	assert RAM(23964) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23964))))  severity failure;
	assert RAM(23965) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(23965))))  severity failure;
	assert RAM(23966) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(23966))))  severity failure;
	assert RAM(23967) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23967))))  severity failure;
	assert RAM(23968) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(23968))))  severity failure;
	assert RAM(23969) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23969))))  severity failure;
	assert RAM(23970) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(23970))))  severity failure;
	assert RAM(23971) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23971))))  severity failure;
	assert RAM(23972) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23972))))  severity failure;
	assert RAM(23973) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(23973))))  severity failure;
	assert RAM(23974) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23974))))  severity failure;
	assert RAM(23975) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(23975))))  severity failure;
	assert RAM(23976) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23976))))  severity failure;
	assert RAM(23977) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(23977))))  severity failure;
	assert RAM(23978) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(23978))))  severity failure;
	assert RAM(23979) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23979))))  severity failure;
	assert RAM(23980) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23980))))  severity failure;
	assert RAM(23981) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23981))))  severity failure;
	assert RAM(23982) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(23982))))  severity failure;
	assert RAM(23983) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23983))))  severity failure;
	assert RAM(23984) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23984))))  severity failure;
	assert RAM(23985) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23985))))  severity failure;
	assert RAM(23986) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(23986))))  severity failure;
	assert RAM(23987) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23987))))  severity failure;
	assert RAM(23988) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(23988))))  severity failure;
	assert RAM(23989) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(23989))))  severity failure;
	assert RAM(23990) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(23990))))  severity failure;
	assert RAM(23991) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(23991))))  severity failure;
	assert RAM(23992) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(23992))))  severity failure;
	assert RAM(23993) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23993))))  severity failure;
	assert RAM(23994) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23994))))  severity failure;
	assert RAM(23995) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23995))))  severity failure;
	assert RAM(23996) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(23996))))  severity failure;
	assert RAM(23997) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23997))))  severity failure;
	assert RAM(23998) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23998))))  severity failure;
	assert RAM(23999) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23999))))  severity failure;
	assert RAM(24000) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24000))))  severity failure;
	assert RAM(24001) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24001))))  severity failure;
	assert RAM(24002) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(24002))))  severity failure;
	assert RAM(24003) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24003))))  severity failure;
	assert RAM(24004) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(24004))))  severity failure;
	assert RAM(24005) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(24005))))  severity failure;
	assert RAM(24006) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(24006))))  severity failure;
	assert RAM(24007) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(24007))))  severity failure;
	assert RAM(24008) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(24008))))  severity failure;
	assert RAM(24009) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24009))))  severity failure;
	assert RAM(24010) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(24010))))  severity failure;
	assert RAM(24011) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(24011))))  severity failure;
	assert RAM(24012) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24012))))  severity failure;
	assert RAM(24013) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(24013))))  severity failure;
	assert RAM(24014) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24014))))  severity failure;
	assert RAM(24015) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24015))))  severity failure;
	assert RAM(24016) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(24016))))  severity failure;
	assert RAM(24017) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24017))))  severity failure;
	assert RAM(24018) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(24018))))  severity failure;
	assert RAM(24019) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24019))))  severity failure;
	assert RAM(24020) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(24020))))  severity failure;
	assert RAM(24021) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(24021))))  severity failure;
	assert RAM(24022) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24022))))  severity failure;
	assert RAM(24023) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(24023))))  severity failure;
	assert RAM(24024) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24024))))  severity failure;
	assert RAM(24025) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(24025))))  severity failure;
	assert RAM(24026) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24026))))  severity failure;
	assert RAM(24027) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(24027))))  severity failure;
	assert RAM(24028) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(24028))))  severity failure;
	assert RAM(24029) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(24029))))  severity failure;
	assert RAM(24030) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24030))))  severity failure;
	assert RAM(24031) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(24031))))  severity failure;
	assert RAM(24032) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24032))))  severity failure;
	assert RAM(24033) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24033))))  severity failure;
	assert RAM(24034) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(24034))))  severity failure;
	assert RAM(24035) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24035))))  severity failure;
	assert RAM(24036) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(24036))))  severity failure;
	assert RAM(24037) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24037))))  severity failure;
	assert RAM(24038) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24038))))  severity failure;
	assert RAM(24039) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24039))))  severity failure;
	assert RAM(24040) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(24040))))  severity failure;
	assert RAM(24041) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(24041))))  severity failure;
	assert RAM(24042) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(24042))))  severity failure;
	assert RAM(24043) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(24043))))  severity failure;
	assert RAM(24044) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(24044))))  severity failure;
	assert RAM(24045) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(24045))))  severity failure;
	assert RAM(24046) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(24046))))  severity failure;
	assert RAM(24047) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(24047))))  severity failure;
	assert RAM(24048) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(24048))))  severity failure;
	assert RAM(24049) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(24049))))  severity failure;
	assert RAM(24050) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(24050))))  severity failure;
	assert RAM(24051) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24051))))  severity failure;
	assert RAM(24052) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(24052))))  severity failure;
	assert RAM(24053) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(24053))))  severity failure;
	assert RAM(24054) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24054))))  severity failure;
	assert RAM(24055) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(24055))))  severity failure;
	assert RAM(24056) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(24056))))  severity failure;
	assert RAM(24057) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(24057))))  severity failure;
	assert RAM(24058) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24058))))  severity failure;
	assert RAM(24059) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(24059))))  severity failure;
	assert RAM(24060) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24060))))  severity failure;
	assert RAM(24061) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24061))))  severity failure;
	assert RAM(24062) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24062))))  severity failure;
	assert RAM(24063) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24063))))  severity failure;
	assert RAM(24064) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24064))))  severity failure;
	assert RAM(24065) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(24065))))  severity failure;
	assert RAM(24066) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(24066))))  severity failure;
	assert RAM(24067) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24067))))  severity failure;
	assert RAM(24068) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24068))))  severity failure;
	assert RAM(24069) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24069))))  severity failure;
	assert RAM(24070) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(24070))))  severity failure;
	assert RAM(24071) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(24071))))  severity failure;
	assert RAM(24072) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(24072))))  severity failure;
	assert RAM(24073) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24073))))  severity failure;
	assert RAM(24074) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(24074))))  severity failure;
	assert RAM(24075) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(24075))))  severity failure;
	assert RAM(24076) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(24076))))  severity failure;
	assert RAM(24077) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(24077))))  severity failure;
	assert RAM(24078) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(24078))))  severity failure;
	assert RAM(24079) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(24079))))  severity failure;
	assert RAM(24080) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(24080))))  severity failure;
	assert RAM(24081) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(24081))))  severity failure;
	assert RAM(24082) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24082))))  severity failure;
	assert RAM(24083) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24083))))  severity failure;
	assert RAM(24084) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24084))))  severity failure;
	assert RAM(24085) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(24085))))  severity failure;
	assert RAM(24086) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24086))))  severity failure;
	assert RAM(24087) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24087))))  severity failure;
	assert RAM(24088) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(24088))))  severity failure;
	assert RAM(24089) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(24089))))  severity failure;
	assert RAM(24090) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(24090))))  severity failure;
	assert RAM(24091) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(24091))))  severity failure;
	assert RAM(24092) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(24092))))  severity failure;
	assert RAM(24093) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(24093))))  severity failure;
	assert RAM(24094) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24094))))  severity failure;
	assert RAM(24095) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24095))))  severity failure;
	assert RAM(24096) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(24096))))  severity failure;
	assert RAM(24097) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24097))))  severity failure;
	assert RAM(24098) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(24098))))  severity failure;
	assert RAM(24099) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24099))))  severity failure;
	assert RAM(24100) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24100))))  severity failure;
	assert RAM(24101) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(24101))))  severity failure;
	assert RAM(24102) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(24102))))  severity failure;
	assert RAM(24103) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24103))))  severity failure;
	assert RAM(24104) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(24104))))  severity failure;
	assert RAM(24105) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(24105))))  severity failure;
	assert RAM(24106) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(24106))))  severity failure;
	assert RAM(24107) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24107))))  severity failure;
	assert RAM(24108) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(24108))))  severity failure;
	assert RAM(24109) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(24109))))  severity failure;
	assert RAM(24110) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(24110))))  severity failure;
	assert RAM(24111) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(24111))))  severity failure;
	assert RAM(24112) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24112))))  severity failure;
	assert RAM(24113) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24113))))  severity failure;
	assert RAM(24114) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(24114))))  severity failure;
	assert RAM(24115) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(24115))))  severity failure;
	assert RAM(24116) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(24116))))  severity failure;
	assert RAM(24117) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24117))))  severity failure;
	assert RAM(24118) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(24118))))  severity failure;
	assert RAM(24119) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(24119))))  severity failure;
	assert RAM(24120) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(24120))))  severity failure;
	assert RAM(24121) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(24121))))  severity failure;
	assert RAM(24122) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(24122))))  severity failure;
	assert RAM(24123) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24123))))  severity failure;
	assert RAM(24124) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(24124))))  severity failure;
	assert RAM(24125) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24125))))  severity failure;
	assert RAM(24126) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24126))))  severity failure;
	assert RAM(24127) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(24127))))  severity failure;
	assert RAM(24128) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(24128))))  severity failure;
	assert RAM(24129) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(24129))))  severity failure;
	assert RAM(24130) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24130))))  severity failure;
	assert RAM(24131) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24131))))  severity failure;
	assert RAM(24132) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24132))))  severity failure;
	assert RAM(24133) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(24133))))  severity failure;
	assert RAM(24134) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24134))))  severity failure;
	assert RAM(24135) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(24135))))  severity failure;
	assert RAM(24136) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(24136))))  severity failure;
	assert RAM(24137) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(24137))))  severity failure;
	assert RAM(24138) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(24138))))  severity failure;
	assert RAM(24139) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24139))))  severity failure;
	assert RAM(24140) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(24140))))  severity failure;
	assert RAM(24141) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(24141))))  severity failure;
	assert RAM(24142) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24142))))  severity failure;
	assert RAM(24143) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(24143))))  severity failure;
	assert RAM(24144) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(24144))))  severity failure;
	assert RAM(24145) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24145))))  severity failure;
	assert RAM(24146) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24146))))  severity failure;
	assert RAM(24147) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(24147))))  severity failure;
	assert RAM(24148) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24148))))  severity failure;
	assert RAM(24149) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(24149))))  severity failure;
	assert RAM(24150) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(24150))))  severity failure;
	assert RAM(24151) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24151))))  severity failure;
	assert RAM(24152) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(24152))))  severity failure;
	assert RAM(24153) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(24153))))  severity failure;
	assert RAM(24154) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(24154))))  severity failure;
	assert RAM(24155) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(24155))))  severity failure;
	assert RAM(24156) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24156))))  severity failure;
	assert RAM(24157) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24157))))  severity failure;
	assert RAM(24158) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24158))))  severity failure;
	assert RAM(24159) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(24159))))  severity failure;
	assert RAM(24160) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24160))))  severity failure;
	assert RAM(24161) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24161))))  severity failure;
	assert RAM(24162) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(24162))))  severity failure;
	assert RAM(24163) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24163))))  severity failure;
	assert RAM(24164) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(24164))))  severity failure;
	assert RAM(24165) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(24165))))  severity failure;
	assert RAM(24166) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24166))))  severity failure;
	assert RAM(24167) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(24167))))  severity failure;
	assert RAM(24168) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(24168))))  severity failure;
	assert RAM(24169) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24169))))  severity failure;
	assert RAM(24170) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24170))))  severity failure;
	assert RAM(24171) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(24171))))  severity failure;
	assert RAM(24172) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24172))))  severity failure;
	assert RAM(24173) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(24173))))  severity failure;
	assert RAM(24174) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(24174))))  severity failure;
	assert RAM(24175) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(24175))))  severity failure;
	assert RAM(24176) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(24176))))  severity failure;
	assert RAM(24177) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(24177))))  severity failure;
	assert RAM(24178) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(24178))))  severity failure;
	assert RAM(24179) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(24179))))  severity failure;
	assert RAM(24180) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24180))))  severity failure;
	assert RAM(24181) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(24181))))  severity failure;
	assert RAM(24182) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(24182))))  severity failure;
	assert RAM(24183) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(24183))))  severity failure;
	assert RAM(24184) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24184))))  severity failure;
	assert RAM(24185) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(24185))))  severity failure;
	assert RAM(24186) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(24186))))  severity failure;
	assert RAM(24187) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(24187))))  severity failure;
	assert RAM(24188) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(24188))))  severity failure;
	assert RAM(24189) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(24189))))  severity failure;
	assert RAM(24190) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24190))))  severity failure;
	assert RAM(24191) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24191))))  severity failure;
	assert RAM(24192) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(24192))))  severity failure;
	assert RAM(24193) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(24193))))  severity failure;
	assert RAM(24194) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(24194))))  severity failure;
	assert RAM(24195) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(24195))))  severity failure;
	assert RAM(24196) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(24196))))  severity failure;
	assert RAM(24197) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(24197))))  severity failure;
	assert RAM(24198) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24198))))  severity failure;
	assert RAM(24199) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24199))))  severity failure;
	assert RAM(24200) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(24200))))  severity failure;
	assert RAM(24201) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24201))))  severity failure;
	assert RAM(24202) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(24202))))  severity failure;
	assert RAM(24203) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24203))))  severity failure;
	assert RAM(24204) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24204))))  severity failure;
	assert RAM(24205) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(24205))))  severity failure;
	assert RAM(24206) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(24206))))  severity failure;
	assert RAM(24207) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24207))))  severity failure;
	assert RAM(24208) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24208))))  severity failure;
	assert RAM(24209) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24209))))  severity failure;
	assert RAM(24210) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(24210))))  severity failure;
	assert RAM(24211) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(24211))))  severity failure;
	assert RAM(24212) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24212))))  severity failure;
	assert RAM(24213) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(24213))))  severity failure;
	assert RAM(24214) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(24214))))  severity failure;
	assert RAM(24215) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(24215))))  severity failure;
	assert RAM(24216) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(24216))))  severity failure;
	assert RAM(24217) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(24217))))  severity failure;
	assert RAM(24218) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(24218))))  severity failure;
	assert RAM(24219) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24219))))  severity failure;
	assert RAM(24220) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24220))))  severity failure;
	assert RAM(24221) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(24221))))  severity failure;
	assert RAM(24222) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(24222))))  severity failure;
	assert RAM(24223) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24223))))  severity failure;
	assert RAM(24224) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24224))))  severity failure;
	assert RAM(24225) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(24225))))  severity failure;
	assert RAM(24226) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(24226))))  severity failure;
	assert RAM(24227) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(24227))))  severity failure;
	assert RAM(24228) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24228))))  severity failure;
	assert RAM(24229) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(24229))))  severity failure;
	assert RAM(24230) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(24230))))  severity failure;
	assert RAM(24231) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(24231))))  severity failure;
	assert RAM(24232) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24232))))  severity failure;
	assert RAM(24233) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24233))))  severity failure;
	assert RAM(24234) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(24234))))  severity failure;
	assert RAM(24235) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24235))))  severity failure;
	assert RAM(24236) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(24236))))  severity failure;
	assert RAM(24237) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24237))))  severity failure;
	assert RAM(24238) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(24238))))  severity failure;
	assert RAM(24239) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(24239))))  severity failure;
	assert RAM(24240) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24240))))  severity failure;
	assert RAM(24241) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(24241))))  severity failure;
	assert RAM(24242) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(24242))))  severity failure;
	assert RAM(24243) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(24243))))  severity failure;
	assert RAM(24244) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(24244))))  severity failure;
	assert RAM(24245) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24245))))  severity failure;
	assert RAM(24246) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(24246))))  severity failure;
	assert RAM(24247) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24247))))  severity failure;
	assert RAM(24248) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(24248))))  severity failure;
	assert RAM(24249) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(24249))))  severity failure;
	assert RAM(24250) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24250))))  severity failure;
	assert RAM(24251) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(24251))))  severity failure;
	assert RAM(24252) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(24252))))  severity failure;
	assert RAM(24253) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(24253))))  severity failure;
	assert RAM(24254) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(24254))))  severity failure;
	assert RAM(24255) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24255))))  severity failure;
	assert RAM(24256) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(24256))))  severity failure;
	assert RAM(24257) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24257))))  severity failure;
	assert RAM(24258) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(24258))))  severity failure;
	assert RAM(24259) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24259))))  severity failure;
	assert RAM(24260) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24260))))  severity failure;
	assert RAM(24261) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(24261))))  severity failure;
	assert RAM(24262) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(24262))))  severity failure;
	assert RAM(24263) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24263))))  severity failure;
	assert RAM(24264) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24264))))  severity failure;
	assert RAM(24265) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24265))))  severity failure;
	assert RAM(24266) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(24266))))  severity failure;
	assert RAM(24267) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(24267))))  severity failure;
	assert RAM(24268) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(24268))))  severity failure;
	assert RAM(24269) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(24269))))  severity failure;
	assert RAM(24270) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24270))))  severity failure;
	assert RAM(24271) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24271))))  severity failure;
	assert RAM(24272) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(24272))))  severity failure;
	assert RAM(24273) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(24273))))  severity failure;
	assert RAM(24274) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(24274))))  severity failure;
	assert RAM(24275) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(24275))))  severity failure;
	assert RAM(24276) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24276))))  severity failure;
	assert RAM(24277) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24277))))  severity failure;
	assert RAM(24278) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(24278))))  severity failure;
	assert RAM(24279) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(24279))))  severity failure;
	assert RAM(24280) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(24280))))  severity failure;
	assert RAM(24281) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(24281))))  severity failure;
	assert RAM(24282) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(24282))))  severity failure;
	assert RAM(24283) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(24283))))  severity failure;
	assert RAM(24284) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(24284))))  severity failure;
	assert RAM(24285) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(24285))))  severity failure;
	assert RAM(24286) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24286))))  severity failure;
	assert RAM(24287) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(24287))))  severity failure;
	assert RAM(24288) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(24288))))  severity failure;
	assert RAM(24289) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24289))))  severity failure;
	assert RAM(24290) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24290))))  severity failure;
	assert RAM(24291) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24291))))  severity failure;
	assert RAM(24292) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(24292))))  severity failure;
	assert RAM(24293) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24293))))  severity failure;
	assert RAM(24294) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(24294))))  severity failure;
	assert RAM(24295) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24295))))  severity failure;
	assert RAM(24296) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(24296))))  severity failure;
	assert RAM(24297) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24297))))  severity failure;
	assert RAM(24298) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(24298))))  severity failure;
	assert RAM(24299) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(24299))))  severity failure;
	assert RAM(24300) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(24300))))  severity failure;
	assert RAM(24301) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(24301))))  severity failure;
	assert RAM(24302) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(24302))))  severity failure;
	assert RAM(24303) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(24303))))  severity failure;
	assert RAM(24304) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24304))))  severity failure;
	assert RAM(24305) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(24305))))  severity failure;
	assert RAM(24306) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(24306))))  severity failure;
	assert RAM(24307) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24307))))  severity failure;
	assert RAM(24308) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24308))))  severity failure;
	assert RAM(24309) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(24309))))  severity failure;
	assert RAM(24310) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24310))))  severity failure;
	assert RAM(24311) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24311))))  severity failure;
	assert RAM(24312) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(24312))))  severity failure;
	assert RAM(24313) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(24313))))  severity failure;
	assert RAM(24314) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24314))))  severity failure;
	assert RAM(24315) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(24315))))  severity failure;
	assert RAM(24316) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24316))))  severity failure;
	assert RAM(24317) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(24317))))  severity failure;
	assert RAM(24318) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(24318))))  severity failure;
	assert RAM(24319) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(24319))))  severity failure;
	assert RAM(24320) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24320))))  severity failure;
	assert RAM(24321) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(24321))))  severity failure;
	assert RAM(24322) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(24322))))  severity failure;
	assert RAM(24323) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24323))))  severity failure;
	assert RAM(24324) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24324))))  severity failure;
	assert RAM(24325) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(24325))))  severity failure;
	assert RAM(24326) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(24326))))  severity failure;
	assert RAM(24327) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24327))))  severity failure;
	assert RAM(24328) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(24328))))  severity failure;
	assert RAM(24329) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(24329))))  severity failure;
	assert RAM(24330) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(24330))))  severity failure;
	assert RAM(24331) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(24331))))  severity failure;
	assert RAM(24332) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(24332))))  severity failure;
	assert RAM(24333) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(24333))))  severity failure;
	assert RAM(24334) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24334))))  severity failure;
	assert RAM(24335) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(24335))))  severity failure;
	assert RAM(24336) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(24336))))  severity failure;
	assert RAM(24337) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24337))))  severity failure;
	assert RAM(24338) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24338))))  severity failure;
	assert RAM(24339) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24339))))  severity failure;
	assert RAM(24340) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24340))))  severity failure;
	assert RAM(24341) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(24341))))  severity failure;
	assert RAM(24342) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(24342))))  severity failure;
	assert RAM(24343) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24343))))  severity failure;
	assert RAM(24344) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(24344))))  severity failure;
	assert RAM(24345) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(24345))))  severity failure;
	assert RAM(24346) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(24346))))  severity failure;
	assert RAM(24347) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24347))))  severity failure;
	assert RAM(24348) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(24348))))  severity failure;
	assert RAM(24349) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(24349))))  severity failure;
	assert RAM(24350) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(24350))))  severity failure;
	assert RAM(24351) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24351))))  severity failure;
	assert RAM(24352) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(24352))))  severity failure;
	assert RAM(24353) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(24353))))  severity failure;
	assert RAM(24354) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(24354))))  severity failure;
	assert RAM(24355) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24355))))  severity failure;
	assert RAM(24356) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24356))))  severity failure;
	assert RAM(24357) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(24357))))  severity failure;
	assert RAM(24358) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24358))))  severity failure;
	assert RAM(24359) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24359))))  severity failure;
	assert RAM(24360) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24360))))  severity failure;
	assert RAM(24361) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24361))))  severity failure;
	assert RAM(24362) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24362))))  severity failure;
	assert RAM(24363) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(24363))))  severity failure;
	assert RAM(24364) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24364))))  severity failure;
	assert RAM(24365) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(24365))))  severity failure;
	assert RAM(24366) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(24366))))  severity failure;
	assert RAM(24367) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24367))))  severity failure;
	assert RAM(24368) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24368))))  severity failure;
	assert RAM(24369) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(24369))))  severity failure;
	assert RAM(24370) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24370))))  severity failure;
	assert RAM(24371) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(24371))))  severity failure;
	assert RAM(24372) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(24372))))  severity failure;
	assert RAM(24373) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(24373))))  severity failure;
	assert RAM(24374) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(24374))))  severity failure;
	assert RAM(24375) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(24375))))  severity failure;
	assert RAM(24376) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24376))))  severity failure;
	assert RAM(24377) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(24377))))  severity failure;
	assert RAM(24378) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24378))))  severity failure;
	assert RAM(24379) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(24379))))  severity failure;
	assert RAM(24380) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(24380))))  severity failure;
	assert RAM(24381) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24381))))  severity failure;
	assert RAM(24382) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(24382))))  severity failure;
	assert RAM(24383) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(24383))))  severity failure;
	assert RAM(24384) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24384))))  severity failure;
	assert RAM(24385) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(24385))))  severity failure;
	assert RAM(24386) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(24386))))  severity failure;
	assert RAM(24387) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(24387))))  severity failure;
	assert RAM(24388) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(24388))))  severity failure;
	assert RAM(24389) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(24389))))  severity failure;
	assert RAM(24390) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24390))))  severity failure;
	assert RAM(24391) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(24391))))  severity failure;
	assert RAM(24392) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(24392))))  severity failure;
	assert RAM(24393) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(24393))))  severity failure;
	assert RAM(24394) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(24394))))  severity failure;
	assert RAM(24395) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(24395))))  severity failure;
	assert RAM(24396) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24396))))  severity failure;
	assert RAM(24397) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24397))))  severity failure;
	assert RAM(24398) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24398))))  severity failure;
	assert RAM(24399) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(24399))))  severity failure;
	assert RAM(24400) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24400))))  severity failure;
	assert RAM(24401) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24401))))  severity failure;
	assert RAM(24402) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(24402))))  severity failure;
	assert RAM(24403) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(24403))))  severity failure;
	assert RAM(24404) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(24404))))  severity failure;
	assert RAM(24405) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24405))))  severity failure;
	assert RAM(24406) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(24406))))  severity failure;
	assert RAM(24407) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24407))))  severity failure;
	assert RAM(24408) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(24408))))  severity failure;
	assert RAM(24409) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(24409))))  severity failure;
	assert RAM(24410) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(24410))))  severity failure;
	assert RAM(24411) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(24411))))  severity failure;
	assert RAM(24412) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24412))))  severity failure;
	assert RAM(24413) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24413))))  severity failure;
	assert RAM(24414) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(24414))))  severity failure;
	assert RAM(24415) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(24415))))  severity failure;
	assert RAM(24416) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(24416))))  severity failure;
	assert RAM(24417) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(24417))))  severity failure;
	assert RAM(24418) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24418))))  severity failure;
	assert RAM(24419) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24419))))  severity failure;
	assert RAM(24420) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24420))))  severity failure;
	assert RAM(24421) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(24421))))  severity failure;
	assert RAM(24422) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(24422))))  severity failure;
	assert RAM(24423) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24423))))  severity failure;
	assert RAM(24424) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24424))))  severity failure;
	assert RAM(24425) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(24425))))  severity failure;
	assert RAM(24426) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(24426))))  severity failure;
	assert RAM(24427) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24427))))  severity failure;
	assert RAM(24428) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24428))))  severity failure;
	assert RAM(24429) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24429))))  severity failure;
	assert RAM(24430) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24430))))  severity failure;
	assert RAM(24431) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(24431))))  severity failure;
	assert RAM(24432) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(24432))))  severity failure;
	assert RAM(24433) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(24433))))  severity failure;
	assert RAM(24434) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(24434))))  severity failure;
	assert RAM(24435) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(24435))))  severity failure;
	assert RAM(24436) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(24436))))  severity failure;
	assert RAM(24437) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(24437))))  severity failure;
	assert RAM(24438) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24438))))  severity failure;
	assert RAM(24439) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(24439))))  severity failure;
	assert RAM(24440) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(24440))))  severity failure;
	assert RAM(24441) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(24441))))  severity failure;
	assert RAM(24442) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24442))))  severity failure;
	assert RAM(24443) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(24443))))  severity failure;
	assert RAM(24444) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24444))))  severity failure;
	assert RAM(24445) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(24445))))  severity failure;
	assert RAM(24446) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24446))))  severity failure;
	assert RAM(24447) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24447))))  severity failure;
	assert RAM(24448) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24448))))  severity failure;
	assert RAM(24449) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(24449))))  severity failure;
	assert RAM(24450) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(24450))))  severity failure;
	assert RAM(24451) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(24451))))  severity failure;
	assert RAM(24452) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24452))))  severity failure;
	assert RAM(24453) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(24453))))  severity failure;
	assert RAM(24454) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(24454))))  severity failure;
	assert RAM(24455) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(24455))))  severity failure;
	assert RAM(24456) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(24456))))  severity failure;
	assert RAM(24457) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(24457))))  severity failure;
	assert RAM(24458) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(24458))))  severity failure;
	assert RAM(24459) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(24459))))  severity failure;
	assert RAM(24460) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(24460))))  severity failure;
	assert RAM(24461) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24461))))  severity failure;
	assert RAM(24462) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24462))))  severity failure;
	assert RAM(24463) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(24463))))  severity failure;
	assert RAM(24464) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(24464))))  severity failure;
	assert RAM(24465) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(24465))))  severity failure;
	assert RAM(24466) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(24466))))  severity failure;
	assert RAM(24467) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(24467))))  severity failure;
	assert RAM(24468) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24468))))  severity failure;
	assert RAM(24469) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(24469))))  severity failure;
	assert RAM(24470) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(24470))))  severity failure;
	assert RAM(24471) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(24471))))  severity failure;
	assert RAM(24472) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(24472))))  severity failure;
	assert RAM(24473) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(24473))))  severity failure;
	assert RAM(24474) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(24474))))  severity failure;
	assert RAM(24475) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24475))))  severity failure;
	assert RAM(24476) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24476))))  severity failure;
	assert RAM(24477) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(24477))))  severity failure;
	assert RAM(24478) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(24478))))  severity failure;
	assert RAM(24479) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(24479))))  severity failure;
	assert RAM(24480) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(24480))))  severity failure;
	assert RAM(24481) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24481))))  severity failure;
	assert RAM(24482) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24482))))  severity failure;
	assert RAM(24483) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(24483))))  severity failure;
	assert RAM(24484) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(24484))))  severity failure;
	assert RAM(24485) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24485))))  severity failure;
	assert RAM(24486) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(24486))))  severity failure;
	assert RAM(24487) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(24487))))  severity failure;
	assert RAM(24488) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(24488))))  severity failure;
	assert RAM(24489) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(24489))))  severity failure;
	assert RAM(24490) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24490))))  severity failure;
	assert RAM(24491) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(24491))))  severity failure;
	assert RAM(24492) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(24492))))  severity failure;
	assert RAM(24493) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(24493))))  severity failure;
	assert RAM(24494) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24494))))  severity failure;
	assert RAM(24495) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24495))))  severity failure;
	assert RAM(24496) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(24496))))  severity failure;
	assert RAM(24497) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(24497))))  severity failure;
	assert RAM(24498) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24498))))  severity failure;
	assert RAM(24499) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(24499))))  severity failure;
	assert RAM(24500) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24500))))  severity failure;
	assert RAM(24501) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24501))))  severity failure;
	assert RAM(24502) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24502))))  severity failure;
	assert RAM(24503) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(24503))))  severity failure;
	assert RAM(24504) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(24504))))  severity failure;
	assert RAM(24505) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(24505))))  severity failure;
	assert RAM(24506) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(24506))))  severity failure;
	assert RAM(24507) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24507))))  severity failure;
	assert RAM(24508) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(24508))))  severity failure;
	assert RAM(24509) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24509))))  severity failure;
	assert RAM(24510) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(24510))))  severity failure;
	assert RAM(24511) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24511))))  severity failure;
	assert RAM(24512) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24512))))  severity failure;
	assert RAM(24513) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(24513))))  severity failure;
	assert RAM(24514) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(24514))))  severity failure;
	assert RAM(24515) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(24515))))  severity failure;
	assert RAM(24516) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24516))))  severity failure;
	assert RAM(24517) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(24517))))  severity failure;
	assert RAM(24518) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(24518))))  severity failure;
	assert RAM(24519) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24519))))  severity failure;
	assert RAM(24520) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(24520))))  severity failure;
	assert RAM(24521) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(24521))))  severity failure;
	assert RAM(24522) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(24522))))  severity failure;
	assert RAM(24523) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(24523))))  severity failure;
	assert RAM(24524) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(24524))))  severity failure;
	assert RAM(24525) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24525))))  severity failure;
	assert RAM(24526) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(24526))))  severity failure;
	assert RAM(24527) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(24527))))  severity failure;
	assert RAM(24528) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(24528))))  severity failure;
	assert RAM(24529) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(24529))))  severity failure;
	assert RAM(24530) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24530))))  severity failure;
	assert RAM(24531) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(24531))))  severity failure;
	assert RAM(24532) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(24532))))  severity failure;
	assert RAM(24533) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(24533))))  severity failure;
	assert RAM(24534) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24534))))  severity failure;
	assert RAM(24535) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(24535))))  severity failure;
	assert RAM(24536) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(24536))))  severity failure;
	assert RAM(24537) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(24537))))  severity failure;
	assert RAM(24538) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(24538))))  severity failure;
	assert RAM(24539) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24539))))  severity failure;
	assert RAM(24540) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(24540))))  severity failure;
	assert RAM(24541) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(24541))))  severity failure;
	assert RAM(24542) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24542))))  severity failure;
	assert RAM(24543) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(24543))))  severity failure;
	assert RAM(24544) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(24544))))  severity failure;
	assert RAM(24545) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(24545))))  severity failure;
	assert RAM(24546) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(24546))))  severity failure;
	assert RAM(24547) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(24547))))  severity failure;
	assert RAM(24548) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24548))))  severity failure;
	assert RAM(24549) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24549))))  severity failure;
	assert RAM(24550) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24550))))  severity failure;
	assert RAM(24551) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(24551))))  severity failure;
	assert RAM(24552) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(24552))))  severity failure;
	assert RAM(24553) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(24553))))  severity failure;
	assert RAM(24554) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(24554))))  severity failure;
	assert RAM(24555) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(24555))))  severity failure;
	assert RAM(24556) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24556))))  severity failure;
	assert RAM(24557) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(24557))))  severity failure;
	assert RAM(24558) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24558))))  severity failure;
	assert RAM(24559) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(24559))))  severity failure;
	assert RAM(24560) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(24560))))  severity failure;
	assert RAM(24561) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24561))))  severity failure;
	assert RAM(24562) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(24562))))  severity failure;
	assert RAM(24563) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(24563))))  severity failure;
	assert RAM(24564) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(24564))))  severity failure;
	assert RAM(24565) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(24565))))  severity failure;
	assert RAM(24566) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24566))))  severity failure;
	assert RAM(24567) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(24567))))  severity failure;
	assert RAM(24568) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(24568))))  severity failure;
	assert RAM(24569) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24569))))  severity failure;
	assert RAM(24570) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(24570))))  severity failure;
	assert RAM(24571) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(24571))))  severity failure;
	assert RAM(24572) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(24572))))  severity failure;
	assert RAM(24573) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(24573))))  severity failure;
	assert RAM(24574) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(24574))))  severity failure;
	assert RAM(24575) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24575))))  severity failure;
	assert RAM(24576) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24576))))  severity failure;
	assert RAM(24577) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(24577))))  severity failure;
	assert RAM(24578) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(24578))))  severity failure;
	assert RAM(24579) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(24579))))  severity failure;
	assert RAM(24580) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(24580))))  severity failure;
	assert RAM(24581) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(24581))))  severity failure;
	assert RAM(24582) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24582))))  severity failure;
	assert RAM(24583) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(24583))))  severity failure;
	assert RAM(24584) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(24584))))  severity failure;
	assert RAM(24585) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(24585))))  severity failure;
	assert RAM(24586) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(24586))))  severity failure;
	assert RAM(24587) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24587))))  severity failure;
	assert RAM(24588) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24588))))  severity failure;
	assert RAM(24589) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24589))))  severity failure;
	assert RAM(24590) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(24590))))  severity failure;
	assert RAM(24591) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(24591))))  severity failure;
	assert RAM(24592) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(24592))))  severity failure;
	assert RAM(24593) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(24593))))  severity failure;
	assert RAM(24594) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(24594))))  severity failure;
	assert RAM(24595) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24595))))  severity failure;
	assert RAM(24596) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(24596))))  severity failure;
	assert RAM(24597) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24597))))  severity failure;
	assert RAM(24598) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(24598))))  severity failure;
	assert RAM(24599) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24599))))  severity failure;
	assert RAM(24600) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24600))))  severity failure;
	assert RAM(24601) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(24601))))  severity failure;
	assert RAM(24602) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(24602))))  severity failure;
	assert RAM(24603) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(24603))))  severity failure;
	assert RAM(24604) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24604))))  severity failure;
	assert RAM(24605) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24605))))  severity failure;
	assert RAM(24606) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(24606))))  severity failure;
	assert RAM(24607) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(24607))))  severity failure;
	assert RAM(24608) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24608))))  severity failure;
	assert RAM(24609) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24609))))  severity failure;
	assert RAM(24610) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24610))))  severity failure;
	assert RAM(24611) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24611))))  severity failure;
	assert RAM(24612) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(24612))))  severity failure;
	assert RAM(24613) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(24613))))  severity failure;
	assert RAM(24614) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(24614))))  severity failure;
	assert RAM(24615) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(24615))))  severity failure;
	assert RAM(24616) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(24616))))  severity failure;
	assert RAM(24617) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24617))))  severity failure;
	assert RAM(24618) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24618))))  severity failure;
	assert RAM(24619) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24619))))  severity failure;
	assert RAM(24620) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24620))))  severity failure;
	assert RAM(24621) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(24621))))  severity failure;
	assert RAM(24622) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(24622))))  severity failure;
	assert RAM(24623) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(24623))))  severity failure;
	assert RAM(24624) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(24624))))  severity failure;
	assert RAM(24625) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(24625))))  severity failure;
	assert RAM(24626) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(24626))))  severity failure;
	assert RAM(24627) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(24627))))  severity failure;
	assert RAM(24628) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24628))))  severity failure;
	assert RAM(24629) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24629))))  severity failure;
	assert RAM(24630) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(24630))))  severity failure;
	assert RAM(24631) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(24631))))  severity failure;
	assert RAM(24632) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24632))))  severity failure;
	assert RAM(24633) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(24633))))  severity failure;
	assert RAM(24634) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(24634))))  severity failure;
	assert RAM(24635) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24635))))  severity failure;
	assert RAM(24636) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(24636))))  severity failure;
	assert RAM(24637) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(24637))))  severity failure;
	assert RAM(24638) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24638))))  severity failure;
	assert RAM(24639) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(24639))))  severity failure;
	assert RAM(24640) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24640))))  severity failure;
	assert RAM(24641) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(24641))))  severity failure;
	assert RAM(24642) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(24642))))  severity failure;
	assert RAM(24643) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24643))))  severity failure;
	assert RAM(24644) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24644))))  severity failure;
	assert RAM(24645) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24645))))  severity failure;
	assert RAM(24646) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24646))))  severity failure;
	assert RAM(24647) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24647))))  severity failure;
	assert RAM(24648) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(24648))))  severity failure;
	assert RAM(24649) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24649))))  severity failure;
	assert RAM(24650) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(24650))))  severity failure;
	assert RAM(24651) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(24651))))  severity failure;
	assert RAM(24652) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(24652))))  severity failure;
	assert RAM(24653) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(24653))))  severity failure;
	assert RAM(24654) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(24654))))  severity failure;
	assert RAM(24655) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(24655))))  severity failure;
	assert RAM(24656) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24656))))  severity failure;
	assert RAM(24657) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(24657))))  severity failure;
	assert RAM(24658) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(24658))))  severity failure;
	assert RAM(24659) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(24659))))  severity failure;
	assert RAM(24660) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(24660))))  severity failure;
	assert RAM(24661) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24661))))  severity failure;
	assert RAM(24662) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(24662))))  severity failure;
	assert RAM(24663) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24663))))  severity failure;
	assert RAM(24664) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(24664))))  severity failure;
	assert RAM(24665) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(24665))))  severity failure;
	assert RAM(24666) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(24666))))  severity failure;
	assert RAM(24667) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24667))))  severity failure;
	assert RAM(24668) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(24668))))  severity failure;
	assert RAM(24669) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24669))))  severity failure;
	assert RAM(24670) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(24670))))  severity failure;
	assert RAM(24671) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(24671))))  severity failure;
	assert RAM(24672) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(24672))))  severity failure;
	assert RAM(24673) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(24673))))  severity failure;
	assert RAM(24674) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(24674))))  severity failure;
	assert RAM(24675) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(24675))))  severity failure;
	assert RAM(24676) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(24676))))  severity failure;
	assert RAM(24677) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(24677))))  severity failure;
	assert RAM(24678) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(24678))))  severity failure;
	assert RAM(24679) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(24679))))  severity failure;
	assert RAM(24680) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(24680))))  severity failure;
	assert RAM(24681) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(24681))))  severity failure;
	assert RAM(24682) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(24682))))  severity failure;
	assert RAM(24683) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(24683))))  severity failure;
	assert RAM(24684) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(24684))))  severity failure;
	assert RAM(24685) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(24685))))  severity failure;
	assert RAM(24686) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(24686))))  severity failure;
	assert RAM(24687) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(24687))))  severity failure;
	assert RAM(24688) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(24688))))  severity failure;
	assert RAM(24689) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(24689))))  severity failure;
	assert RAM(24690) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(24690))))  severity failure;
	assert RAM(24691) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(24691))))  severity failure;
	assert RAM(24692) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(24692))))  severity failure;
	assert RAM(24693) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(24693))))  severity failure;
	assert RAM(24694) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24694))))  severity failure;
	assert RAM(24695) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(24695))))  severity failure;
	assert RAM(24696) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24696))))  severity failure;
	assert RAM(24697) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(24697))))  severity failure;
	assert RAM(24698) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(24698))))  severity failure;
	assert RAM(24699) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24699))))  severity failure;
	assert RAM(24700) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(24700))))  severity failure;
	assert RAM(24701) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(24701))))  severity failure;
	assert RAM(24702) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(24702))))  severity failure;
	assert RAM(24703) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24703))))  severity failure;
	assert RAM(24704) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24704))))  severity failure;
	assert RAM(24705) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(24705))))  severity failure;
	assert RAM(24706) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(24706))))  severity failure;
	assert RAM(24707) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24707))))  severity failure;
	assert RAM(24708) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24708))))  severity failure;
	assert RAM(24709) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(24709))))  severity failure;
	assert RAM(24710) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(24710))))  severity failure;
	assert RAM(24711) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(24711))))  severity failure;
	assert RAM(24712) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(24712))))  severity failure;
	assert RAM(24713) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(24713))))  severity failure;
	assert RAM(24714) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(24714))))  severity failure;
	assert RAM(24715) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(24715))))  severity failure;
	assert RAM(24716) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24716))))  severity failure;
	assert RAM(24717) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(24717))))  severity failure;
	assert RAM(24718) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(24718))))  severity failure;
	assert RAM(24719) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24719))))  severity failure;
	assert RAM(24720) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(24720))))  severity failure;
	assert RAM(24721) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24721))))  severity failure;
	assert RAM(24722) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24722))))  severity failure;
	assert RAM(24723) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24723))))  severity failure;
	assert RAM(24724) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24724))))  severity failure;
	assert RAM(24725) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(24725))))  severity failure;
	assert RAM(24726) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(24726))))  severity failure;
	assert RAM(24727) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24727))))  severity failure;
	assert RAM(24728) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(24728))))  severity failure;
	assert RAM(24729) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(24729))))  severity failure;
	assert RAM(24730) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(24730))))  severity failure;
	assert RAM(24731) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(24731))))  severity failure;
	assert RAM(24732) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(24732))))  severity failure;
	assert RAM(24733) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24733))))  severity failure;
	assert RAM(24734) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(24734))))  severity failure;
	assert RAM(24735) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24735))))  severity failure;
	assert RAM(24736) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(24736))))  severity failure;
	assert RAM(24737) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24737))))  severity failure;
	assert RAM(24738) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24738))))  severity failure;
	assert RAM(24739) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(24739))))  severity failure;
	assert RAM(24740) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(24740))))  severity failure;
	assert RAM(24741) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24741))))  severity failure;
	assert RAM(24742) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(24742))))  severity failure;
	assert RAM(24743) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(24743))))  severity failure;
	assert RAM(24744) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(24744))))  severity failure;
	assert RAM(24745) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24745))))  severity failure;
	assert RAM(24746) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(24746))))  severity failure;
	assert RAM(24747) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(24747))))  severity failure;
	assert RAM(24748) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(24748))))  severity failure;
	assert RAM(24749) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(24749))))  severity failure;
	assert RAM(24750) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24750))))  severity failure;
	assert RAM(24751) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(24751))))  severity failure;
	assert RAM(24752) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24752))))  severity failure;
	assert RAM(24753) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24753))))  severity failure;
	assert RAM(24754) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24754))))  severity failure;
	assert RAM(24755) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(24755))))  severity failure;
	assert RAM(24756) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(24756))))  severity failure;
	assert RAM(24757) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(24757))))  severity failure;
	assert RAM(24758) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(24758))))  severity failure;
	assert RAM(24759) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(24759))))  severity failure;
	assert RAM(24760) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(24760))))  severity failure;
	assert RAM(24761) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24761))))  severity failure;
	assert RAM(24762) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(24762))))  severity failure;
	assert RAM(24763) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(24763))))  severity failure;
	assert RAM(24764) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24764))))  severity failure;
	assert RAM(24765) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(24765))))  severity failure;
	assert RAM(24766) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24766))))  severity failure;
	assert RAM(24767) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(24767))))  severity failure;
	assert RAM(24768) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(24768))))  severity failure;
	assert RAM(24769) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(24769))))  severity failure;
	assert RAM(24770) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24770))))  severity failure;
	assert RAM(24771) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(24771))))  severity failure;
	assert RAM(24772) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(24772))))  severity failure;
	assert RAM(24773) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(24773))))  severity failure;
	assert RAM(24774) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(24774))))  severity failure;
	assert RAM(24775) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(24775))))  severity failure;
	assert RAM(24776) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24776))))  severity failure;
	assert RAM(24777) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24777))))  severity failure;
	assert RAM(24778) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24778))))  severity failure;
	assert RAM(24779) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(24779))))  severity failure;
	assert RAM(24780) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(24780))))  severity failure;
	assert RAM(24781) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(24781))))  severity failure;
	assert RAM(24782) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(24782))))  severity failure;
	assert RAM(24783) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(24783))))  severity failure;
	assert RAM(24784) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(24784))))  severity failure;
	assert RAM(24785) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24785))))  severity failure;
	assert RAM(24786) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(24786))))  severity failure;
	assert RAM(24787) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(24787))))  severity failure;
	assert RAM(24788) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(24788))))  severity failure;
	assert RAM(24789) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(24789))))  severity failure;
	assert RAM(24790) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(24790))))  severity failure;
	assert RAM(24791) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(24791))))  severity failure;
	assert RAM(24792) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24792))))  severity failure;
	assert RAM(24793) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24793))))  severity failure;
	assert RAM(24794) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(24794))))  severity failure;
	assert RAM(24795) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(24795))))  severity failure;
	assert RAM(24796) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(24796))))  severity failure;
	assert RAM(24797) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(24797))))  severity failure;
	assert RAM(24798) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(24798))))  severity failure;
	assert RAM(24799) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24799))))  severity failure;
	assert RAM(24800) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(24800))))  severity failure;
	assert RAM(24801) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(24801))))  severity failure;
	assert RAM(24802) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(24802))))  severity failure;
	assert RAM(24803) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(24803))))  severity failure;
	assert RAM(24804) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(24804))))  severity failure;
	assert RAM(24805) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(24805))))  severity failure;
	assert RAM(24806) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(24806))))  severity failure;
	assert RAM(24807) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(24807))))  severity failure;
	assert RAM(24808) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(24808))))  severity failure;
	assert RAM(24809) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(24809))))  severity failure;
	assert RAM(24810) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(24810))))  severity failure;
	assert RAM(24811) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(24811))))  severity failure;
	assert RAM(24812) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(24812))))  severity failure;
	assert RAM(24813) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24813))))  severity failure;
	assert RAM(24814) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24814))))  severity failure;
	assert RAM(24815) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24815))))  severity failure;
	assert RAM(24816) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24816))))  severity failure;
	assert RAM(24817) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(24817))))  severity failure;
	assert RAM(24818) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(24818))))  severity failure;
	assert RAM(24819) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(24819))))  severity failure;
	assert RAM(24820) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(24820))))  severity failure;
	assert RAM(24821) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(24821))))  severity failure;
	assert RAM(24822) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(24822))))  severity failure;
	assert RAM(24823) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24823))))  severity failure;
	assert RAM(24824) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(24824))))  severity failure;
	assert RAM(24825) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(24825))))  severity failure;
	assert RAM(24826) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(24826))))  severity failure;
	assert RAM(24827) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(24827))))  severity failure;
	assert RAM(24828) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24828))))  severity failure;
	assert RAM(24829) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(24829))))  severity failure;
	assert RAM(24830) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24830))))  severity failure;
	assert RAM(24831) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24831))))  severity failure;
	assert RAM(24832) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24832))))  severity failure;
	assert RAM(24833) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(24833))))  severity failure;
	assert RAM(24834) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24834))))  severity failure;
	assert RAM(24835) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24835))))  severity failure;
	assert RAM(24836) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24836))))  severity failure;
	assert RAM(24837) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(24837))))  severity failure;
	assert RAM(24838) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24838))))  severity failure;
	assert RAM(24839) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(24839))))  severity failure;
	assert RAM(24840) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24840))))  severity failure;
	assert RAM(24841) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24841))))  severity failure;
	assert RAM(24842) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(24842))))  severity failure;
	assert RAM(24843) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(24843))))  severity failure;
	assert RAM(24844) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(24844))))  severity failure;
	assert RAM(24845) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(24845))))  severity failure;
	assert RAM(24846) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24846))))  severity failure;
	assert RAM(24847) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(24847))))  severity failure;
	assert RAM(24848) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(24848))))  severity failure;
	assert RAM(24849) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(24849))))  severity failure;
	assert RAM(24850) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24850))))  severity failure;
	assert RAM(24851) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(24851))))  severity failure;
	assert RAM(24852) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(24852))))  severity failure;
	assert RAM(24853) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(24853))))  severity failure;
	assert RAM(24854) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(24854))))  severity failure;
	assert RAM(24855) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24855))))  severity failure;
	assert RAM(24856) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(24856))))  severity failure;
	assert RAM(24857) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(24857))))  severity failure;
	assert RAM(24858) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24858))))  severity failure;
	assert RAM(24859) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(24859))))  severity failure;
	assert RAM(24860) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(24860))))  severity failure;
	assert RAM(24861) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24861))))  severity failure;
	assert RAM(24862) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(24862))))  severity failure;
	assert RAM(24863) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(24863))))  severity failure;
	assert RAM(24864) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(24864))))  severity failure;
	assert RAM(24865) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(24865))))  severity failure;
	assert RAM(24866) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(24866))))  severity failure;
	assert RAM(24867) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(24867))))  severity failure;
	assert RAM(24868) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(24868))))  severity failure;
	assert RAM(24869) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(24869))))  severity failure;
	assert RAM(24870) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(24870))))  severity failure;
	assert RAM(24871) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(24871))))  severity failure;
	assert RAM(24872) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24872))))  severity failure;
	assert RAM(24873) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(24873))))  severity failure;
	assert RAM(24874) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24874))))  severity failure;
	assert RAM(24875) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(24875))))  severity failure;
	assert RAM(24876) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(24876))))  severity failure;
	assert RAM(24877) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(24877))))  severity failure;
	assert RAM(24878) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(24878))))  severity failure;
	assert RAM(24879) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(24879))))  severity failure;
	assert RAM(24880) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(24880))))  severity failure;
	assert RAM(24881) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(24881))))  severity failure;
	assert RAM(24882) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(24882))))  severity failure;
	assert RAM(24883) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(24883))))  severity failure;
	assert RAM(24884) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(24884))))  severity failure;
	assert RAM(24885) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(24885))))  severity failure;
	assert RAM(24886) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(24886))))  severity failure;
	assert RAM(24887) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24887))))  severity failure;
	assert RAM(24888) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(24888))))  severity failure;
	assert RAM(24889) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(24889))))  severity failure;
	assert RAM(24890) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24890))))  severity failure;
	assert RAM(24891) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(24891))))  severity failure;
	assert RAM(24892) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(24892))))  severity failure;
	assert RAM(24893) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(24893))))  severity failure;
	assert RAM(24894) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(24894))))  severity failure;
	assert RAM(24895) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(24895))))  severity failure;
	assert RAM(24896) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(24896))))  severity failure;
	assert RAM(24897) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(24897))))  severity failure;
	assert RAM(24898) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24898))))  severity failure;
	assert RAM(24899) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24899))))  severity failure;
	assert RAM(24900) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(24900))))  severity failure;
	assert RAM(24901) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24901))))  severity failure;
	assert RAM(24902) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(24902))))  severity failure;
	assert RAM(24903) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(24903))))  severity failure;
	assert RAM(24904) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(24904))))  severity failure;
	assert RAM(24905) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(24905))))  severity failure;
	assert RAM(24906) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24906))))  severity failure;
	assert RAM(24907) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(24907))))  severity failure;
	assert RAM(24908) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(24908))))  severity failure;
	assert RAM(24909) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24909))))  severity failure;
	assert RAM(24910) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(24910))))  severity failure;
	assert RAM(24911) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(24911))))  severity failure;
	assert RAM(24912) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(24912))))  severity failure;
	assert RAM(24913) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(24913))))  severity failure;
	assert RAM(24914) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(24914))))  severity failure;
	assert RAM(24915) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24915))))  severity failure;
	assert RAM(24916) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(24916))))  severity failure;
	assert RAM(24917) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(24917))))  severity failure;
	assert RAM(24918) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(24918))))  severity failure;
	assert RAM(24919) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24919))))  severity failure;
	assert RAM(24920) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(24920))))  severity failure;
	assert RAM(24921) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(24921))))  severity failure;
	assert RAM(24922) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(24922))))  severity failure;
	assert RAM(24923) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(24923))))  severity failure;
	assert RAM(24924) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(24924))))  severity failure;
	assert RAM(24925) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(24925))))  severity failure;
	assert RAM(24926) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24926))))  severity failure;
	assert RAM(24927) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(24927))))  severity failure;
	assert RAM(24928) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(24928))))  severity failure;
	assert RAM(24929) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(24929))))  severity failure;
	assert RAM(24930) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(24930))))  severity failure;
	assert RAM(24931) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(24931))))  severity failure;
	assert RAM(24932) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(24932))))  severity failure;
	assert RAM(24933) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(24933))))  severity failure;
	assert RAM(24934) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24934))))  severity failure;
	assert RAM(24935) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(24935))))  severity failure;
	assert RAM(24936) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(24936))))  severity failure;
	assert RAM(24937) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(24937))))  severity failure;
	assert RAM(24938) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(24938))))  severity failure;
	assert RAM(24939) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(24939))))  severity failure;
	assert RAM(24940) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24940))))  severity failure;
	assert RAM(24941) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(24941))))  severity failure;
	assert RAM(24942) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(24942))))  severity failure;
	assert RAM(24943) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(24943))))  severity failure;
	assert RAM(24944) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(24944))))  severity failure;
	assert RAM(24945) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(24945))))  severity failure;
	assert RAM(24946) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24946))))  severity failure;
	assert RAM(24947) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(24947))))  severity failure;
	assert RAM(24948) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(24948))))  severity failure;
	assert RAM(24949) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(24949))))  severity failure;
	assert RAM(24950) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(24950))))  severity failure;
	assert RAM(24951) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(24951))))  severity failure;
	assert RAM(24952) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(24952))))  severity failure;
	assert RAM(24953) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(24953))))  severity failure;
	assert RAM(24954) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(24954))))  severity failure;
	assert RAM(24955) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(24955))))  severity failure;
	assert RAM(24956) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(24956))))  severity failure;
	assert RAM(24957) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(24957))))  severity failure;
	assert RAM(24958) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(24958))))  severity failure;
	assert RAM(24959) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(24959))))  severity failure;
	assert RAM(24960) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(24960))))  severity failure;
	assert RAM(24961) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(24961))))  severity failure;
	assert RAM(24962) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(24962))))  severity failure;
	assert RAM(24963) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(24963))))  severity failure;
	assert RAM(24964) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(24964))))  severity failure;
	assert RAM(24965) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(24965))))  severity failure;
	assert RAM(24966) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(24966))))  severity failure;
	assert RAM(24967) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(24967))))  severity failure;
	assert RAM(24968) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(24968))))  severity failure;
	assert RAM(24969) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(24969))))  severity failure;
	assert RAM(24970) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(24970))))  severity failure;
	assert RAM(24971) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(24971))))  severity failure;
	assert RAM(24972) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(24972))))  severity failure;
	assert RAM(24973) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(24973))))  severity failure;
	assert RAM(24974) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(24974))))  severity failure;
	assert RAM(24975) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(24975))))  severity failure;
	assert RAM(24976) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(24976))))  severity failure;
	assert RAM(24977) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(24977))))  severity failure;
	assert RAM(24978) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24978))))  severity failure;
	assert RAM(24979) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(24979))))  severity failure;
	assert RAM(24980) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(24980))))  severity failure;
	assert RAM(24981) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(24981))))  severity failure;
	assert RAM(24982) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(24982))))  severity failure;
	assert RAM(24983) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(24983))))  severity failure;
	assert RAM(24984) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(24984))))  severity failure;
	assert RAM(24985) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(24985))))  severity failure;
	assert RAM(24986) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(24986))))  severity failure;
	assert RAM(24987) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(24987))))  severity failure;
	assert RAM(24988) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(24988))))  severity failure;
	assert RAM(24989) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(24989))))  severity failure;
	assert RAM(24990) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(24990))))  severity failure;
	assert RAM(24991) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(24991))))  severity failure;
	assert RAM(24992) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(24992))))  severity failure;
	assert RAM(24993) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(24993))))  severity failure;
	assert RAM(24994) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(24994))))  severity failure;
	assert RAM(24995) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(24995))))  severity failure;
	assert RAM(24996) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(24996))))  severity failure;
	assert RAM(24997) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(24997))))  severity failure;
	assert RAM(24998) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(24998))))  severity failure;
	assert RAM(24999) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(24999))))  severity failure;
	assert RAM(25000) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(25000))))  severity failure;
	assert RAM(25001) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25001))))  severity failure;
	assert RAM(25002) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25002))))  severity failure;
	assert RAM(25003) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(25003))))  severity failure;
	assert RAM(25004) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(25004))))  severity failure;
	assert RAM(25005) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(25005))))  severity failure;
	assert RAM(25006) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25006))))  severity failure;
	assert RAM(25007) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(25007))))  severity failure;
	assert RAM(25008) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(25008))))  severity failure;
	assert RAM(25009) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(25009))))  severity failure;
	assert RAM(25010) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25010))))  severity failure;
	assert RAM(25011) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(25011))))  severity failure;
	assert RAM(25012) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(25012))))  severity failure;
	assert RAM(25013) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(25013))))  severity failure;
	assert RAM(25014) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(25014))))  severity failure;
	assert RAM(25015) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(25015))))  severity failure;
	assert RAM(25016) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(25016))))  severity failure;
	assert RAM(25017) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(25017))))  severity failure;
	assert RAM(25018) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(25018))))  severity failure;
	assert RAM(25019) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25019))))  severity failure;
	assert RAM(25020) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(25020))))  severity failure;
	assert RAM(25021) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(25021))))  severity failure;
	assert RAM(25022) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(25022))))  severity failure;
	assert RAM(25023) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(25023))))  severity failure;
	assert RAM(25024) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25024))))  severity failure;
	assert RAM(25025) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25025))))  severity failure;
	assert RAM(25026) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(25026))))  severity failure;
	assert RAM(25027) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(25027))))  severity failure;
	assert RAM(25028) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(25028))))  severity failure;
	assert RAM(25029) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(25029))))  severity failure;
	assert RAM(25030) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25030))))  severity failure;
	assert RAM(25031) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(25031))))  severity failure;
	assert RAM(25032) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(25032))))  severity failure;
	assert RAM(25033) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25033))))  severity failure;
	assert RAM(25034) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(25034))))  severity failure;
	assert RAM(25035) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(25035))))  severity failure;
	assert RAM(25036) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(25036))))  severity failure;
	assert RAM(25037) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25037))))  severity failure;
	assert RAM(25038) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(25038))))  severity failure;
	assert RAM(25039) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(25039))))  severity failure;
	assert RAM(25040) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(25040))))  severity failure;
	assert RAM(25041) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25041))))  severity failure;
	assert RAM(25042) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(25042))))  severity failure;
	assert RAM(25043) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(25043))))  severity failure;
	assert RAM(25044) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(25044))))  severity failure;
	assert RAM(25045) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(25045))))  severity failure;
	assert RAM(25046) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(25046))))  severity failure;
	assert RAM(25047) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(25047))))  severity failure;
	assert RAM(25048) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(25048))))  severity failure;
	assert RAM(25049) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(25049))))  severity failure;
	assert RAM(25050) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25050))))  severity failure;
	assert RAM(25051) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25051))))  severity failure;
	assert RAM(25052) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25052))))  severity failure;
	assert RAM(25053) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(25053))))  severity failure;
	assert RAM(25054) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25054))))  severity failure;
	assert RAM(25055) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(25055))))  severity failure;
	assert RAM(25056) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(25056))))  severity failure;
	assert RAM(25057) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25057))))  severity failure;
	assert RAM(25058) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(25058))))  severity failure;
	assert RAM(25059) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(25059))))  severity failure;
	assert RAM(25060) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(25060))))  severity failure;
	assert RAM(25061) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25061))))  severity failure;
	assert RAM(25062) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25062))))  severity failure;
	assert RAM(25063) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25063))))  severity failure;
	assert RAM(25064) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(25064))))  severity failure;
	assert RAM(25065) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(25065))))  severity failure;
	assert RAM(25066) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(25066))))  severity failure;
	assert RAM(25067) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25067))))  severity failure;
	assert RAM(25068) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25068))))  severity failure;
	assert RAM(25069) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(25069))))  severity failure;
	assert RAM(25070) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(25070))))  severity failure;
	assert RAM(25071) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25071))))  severity failure;
	assert RAM(25072) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(25072))))  severity failure;
	assert RAM(25073) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25073))))  severity failure;
	assert RAM(25074) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(25074))))  severity failure;
	assert RAM(25075) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(25075))))  severity failure;
	assert RAM(25076) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(25076))))  severity failure;
	assert RAM(25077) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(25077))))  severity failure;
	assert RAM(25078) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(25078))))  severity failure;
	assert RAM(25079) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(25079))))  severity failure;
	assert RAM(25080) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(25080))))  severity failure;
	assert RAM(25081) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(25081))))  severity failure;
	assert RAM(25082) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(25082))))  severity failure;
	assert RAM(25083) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25083))))  severity failure;
	assert RAM(25084) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25084))))  severity failure;
	assert RAM(25085) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25085))))  severity failure;
	assert RAM(25086) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25086))))  severity failure;
	assert RAM(25087) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(25087))))  severity failure;
	assert RAM(25088) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25088))))  severity failure;
	assert RAM(25089) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(25089))))  severity failure;
	assert RAM(25090) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(25090))))  severity failure;
	assert RAM(25091) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(25091))))  severity failure;
	assert RAM(25092) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25092))))  severity failure;
	assert RAM(25093) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25093))))  severity failure;
	assert RAM(25094) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(25094))))  severity failure;
	assert RAM(25095) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25095))))  severity failure;
	assert RAM(25096) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25096))))  severity failure;
	assert RAM(25097) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25097))))  severity failure;
	assert RAM(25098) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25098))))  severity failure;
	assert RAM(25099) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25099))))  severity failure;
	assert RAM(25100) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(25100))))  severity failure;
	assert RAM(25101) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25101))))  severity failure;
	assert RAM(25102) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(25102))))  severity failure;
	assert RAM(25103) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(25103))))  severity failure;
	assert RAM(25104) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25104))))  severity failure;
	assert RAM(25105) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(25105))))  severity failure;
	assert RAM(25106) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25106))))  severity failure;
	assert RAM(25107) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25107))))  severity failure;
	assert RAM(25108) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(25108))))  severity failure;
	assert RAM(25109) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25109))))  severity failure;
	assert RAM(25110) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(25110))))  severity failure;
	assert RAM(25111) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(25111))))  severity failure;
	assert RAM(25112) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(25112))))  severity failure;
	assert RAM(25113) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(25113))))  severity failure;
	assert RAM(25114) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25114))))  severity failure;
	assert RAM(25115) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(25115))))  severity failure;
	assert RAM(25116) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(25116))))  severity failure;
	assert RAM(25117) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(25117))))  severity failure;
	assert RAM(25118) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25118))))  severity failure;
	assert RAM(25119) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(25119))))  severity failure;
	assert RAM(25120) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25120))))  severity failure;
	assert RAM(25121) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(25121))))  severity failure;
	assert RAM(25122) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(25122))))  severity failure;
	assert RAM(25123) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25123))))  severity failure;
	assert RAM(25124) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(25124))))  severity failure;
	assert RAM(25125) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(25125))))  severity failure;
	assert RAM(25126) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(25126))))  severity failure;
	assert RAM(25127) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(25127))))  severity failure;
	assert RAM(25128) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(25128))))  severity failure;
	assert RAM(25129) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(25129))))  severity failure;
	assert RAM(25130) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(25130))))  severity failure;
	assert RAM(25131) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25131))))  severity failure;
	assert RAM(25132) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25132))))  severity failure;
	assert RAM(25133) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(25133))))  severity failure;
	assert RAM(25134) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(25134))))  severity failure;
	assert RAM(25135) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(25135))))  severity failure;
	assert RAM(25136) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(25136))))  severity failure;
	assert RAM(25137) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25137))))  severity failure;
	assert RAM(25138) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(25138))))  severity failure;
	assert RAM(25139) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(25139))))  severity failure;
	assert RAM(25140) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25140))))  severity failure;
	assert RAM(25141) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25141))))  severity failure;
	assert RAM(25142) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(25142))))  severity failure;
	assert RAM(25143) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25143))))  severity failure;
	assert RAM(25144) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(25144))))  severity failure;
	assert RAM(25145) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25145))))  severity failure;
	assert RAM(25146) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(25146))))  severity failure;
	assert RAM(25147) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(25147))))  severity failure;
	assert RAM(25148) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(25148))))  severity failure;
	assert RAM(25149) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(25149))))  severity failure;
	assert RAM(25150) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25150))))  severity failure;
	assert RAM(25151) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(25151))))  severity failure;
	assert RAM(25152) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(25152))))  severity failure;
	assert RAM(25153) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(25153))))  severity failure;
	assert RAM(25154) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(25154))))  severity failure;
	assert RAM(25155) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(25155))))  severity failure;
	assert RAM(25156) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25156))))  severity failure;
	assert RAM(25157) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(25157))))  severity failure;
	assert RAM(25158) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(25158))))  severity failure;
	assert RAM(25159) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(25159))))  severity failure;
	assert RAM(25160) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(25160))))  severity failure;
	assert RAM(25161) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(25161))))  severity failure;
	assert RAM(25162) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25162))))  severity failure;
	assert RAM(25163) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25163))))  severity failure;
	assert RAM(25164) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(25164))))  severity failure;
	assert RAM(25165) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(25165))))  severity failure;
	assert RAM(25166) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(25166))))  severity failure;
	assert RAM(25167) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(25167))))  severity failure;
	assert RAM(25168) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(25168))))  severity failure;
	assert RAM(25169) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25169))))  severity failure;
	assert RAM(25170) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25170))))  severity failure;
	assert RAM(25171) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25171))))  severity failure;
	assert RAM(25172) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(25172))))  severity failure;
	assert RAM(25173) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(25173))))  severity failure;
	assert RAM(25174) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(25174))))  severity failure;
	assert RAM(25175) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25175))))  severity failure;
	assert RAM(25176) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(25176))))  severity failure;
	assert RAM(25177) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(25177))))  severity failure;
	assert RAM(25178) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25178))))  severity failure;
	assert RAM(25179) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(25179))))  severity failure;
	assert RAM(25180) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(25180))))  severity failure;
	assert RAM(25181) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(25181))))  severity failure;
	assert RAM(25182) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(25182))))  severity failure;
	assert RAM(25183) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(25183))))  severity failure;
	assert RAM(25184) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(25184))))  severity failure;
	assert RAM(25185) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25185))))  severity failure;
	assert RAM(25186) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(25186))))  severity failure;
	assert RAM(25187) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(25187))))  severity failure;
	assert RAM(25188) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(25188))))  severity failure;
	assert RAM(25189) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(25189))))  severity failure;
	assert RAM(25190) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25190))))  severity failure;
	assert RAM(25191) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(25191))))  severity failure;
	assert RAM(25192) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(25192))))  severity failure;
	assert RAM(25193) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(25193))))  severity failure;
	assert RAM(25194) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(25194))))  severity failure;
	assert RAM(25195) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25195))))  severity failure;
	assert RAM(25196) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25196))))  severity failure;
	assert RAM(25197) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(25197))))  severity failure;
	assert RAM(25198) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25198))))  severity failure;
	assert RAM(25199) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25199))))  severity failure;
	assert RAM(25200) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(25200))))  severity failure;
	assert RAM(25201) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(25201))))  severity failure;
	assert RAM(25202) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25202))))  severity failure;
	assert RAM(25203) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(25203))))  severity failure;
	assert RAM(25204) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25204))))  severity failure;
	assert RAM(25205) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(25205))))  severity failure;
	assert RAM(25206) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25206))))  severity failure;
	assert RAM(25207) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25207))))  severity failure;
	assert RAM(25208) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25208))))  severity failure;
	assert RAM(25209) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25209))))  severity failure;
	assert RAM(25210) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(25210))))  severity failure;
	assert RAM(25211) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(25211))))  severity failure;
	assert RAM(25212) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(25212))))  severity failure;
	assert RAM(25213) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(25213))))  severity failure;
	assert RAM(25214) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(25214))))  severity failure;
	assert RAM(25215) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25215))))  severity failure;
	assert RAM(25216) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(25216))))  severity failure;
	assert RAM(25217) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(25217))))  severity failure;
	assert RAM(25218) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(25218))))  severity failure;
	assert RAM(25219) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(25219))))  severity failure;
	assert RAM(25220) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(25220))))  severity failure;
	assert RAM(25221) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25221))))  severity failure;
	assert RAM(25222) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(25222))))  severity failure;
	assert RAM(25223) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(25223))))  severity failure;
	assert RAM(25224) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25224))))  severity failure;
	assert RAM(25225) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(25225))))  severity failure;
	assert RAM(25226) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(25226))))  severity failure;
	assert RAM(25227) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(25227))))  severity failure;
	assert RAM(25228) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25228))))  severity failure;
	assert RAM(25229) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(25229))))  severity failure;
	assert RAM(25230) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(25230))))  severity failure;
	assert RAM(25231) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25231))))  severity failure;
	assert RAM(25232) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(25232))))  severity failure;
	assert RAM(25233) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25233))))  severity failure;
	assert RAM(25234) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(25234))))  severity failure;
	assert RAM(25235) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(25235))))  severity failure;
	assert RAM(25236) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(25236))))  severity failure;
	assert RAM(25237) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(25237))))  severity failure;
	assert RAM(25238) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(25238))))  severity failure;
	assert RAM(25239) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(25239))))  severity failure;
	assert RAM(25240) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(25240))))  severity failure;
	assert RAM(25241) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(25241))))  severity failure;
	assert RAM(25242) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(25242))))  severity failure;
	assert RAM(25243) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(25243))))  severity failure;
	assert RAM(25244) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(25244))))  severity failure;
	assert RAM(25245) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(25245))))  severity failure;
	assert RAM(25246) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25246))))  severity failure;
	assert RAM(25247) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(25247))))  severity failure;
	assert RAM(25248) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(25248))))  severity failure;
	assert RAM(25249) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(25249))))  severity failure;
	assert RAM(25250) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25250))))  severity failure;
	assert RAM(25251) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25251))))  severity failure;
	assert RAM(25252) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25252))))  severity failure;
	assert RAM(25253) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(25253))))  severity failure;
	assert RAM(25254) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(25254))))  severity failure;
	assert RAM(25255) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25255))))  severity failure;
	assert RAM(25256) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25256))))  severity failure;
	assert RAM(25257) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25257))))  severity failure;
	assert RAM(25258) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(25258))))  severity failure;
	assert RAM(25259) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(25259))))  severity failure;
	assert RAM(25260) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25260))))  severity failure;
	assert RAM(25261) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(25261))))  severity failure;
	assert RAM(25262) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(25262))))  severity failure;
	assert RAM(25263) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(25263))))  severity failure;
	assert RAM(25264) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(25264))))  severity failure;
	assert RAM(25265) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(25265))))  severity failure;
	assert RAM(25266) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(25266))))  severity failure;
	assert RAM(25267) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25267))))  severity failure;
	assert RAM(25268) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25268))))  severity failure;
	assert RAM(25269) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25269))))  severity failure;
	assert RAM(25270) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25270))))  severity failure;
	assert RAM(25271) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(25271))))  severity failure;
	assert RAM(25272) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(25272))))  severity failure;
	assert RAM(25273) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(25273))))  severity failure;
	assert RAM(25274) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25274))))  severity failure;
	assert RAM(25275) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(25275))))  severity failure;
	assert RAM(25276) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(25276))))  severity failure;
	assert RAM(25277) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(25277))))  severity failure;
	assert RAM(25278) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(25278))))  severity failure;
	assert RAM(25279) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(25279))))  severity failure;
	assert RAM(25280) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(25280))))  severity failure;
	assert RAM(25281) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(25281))))  severity failure;
	assert RAM(25282) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25282))))  severity failure;
	assert RAM(25283) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(25283))))  severity failure;
	assert RAM(25284) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(25284))))  severity failure;
	assert RAM(25285) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(25285))))  severity failure;
	assert RAM(25286) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(25286))))  severity failure;
	assert RAM(25287) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25287))))  severity failure;
	assert RAM(25288) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(25288))))  severity failure;
	assert RAM(25289) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(25289))))  severity failure;
	assert RAM(25290) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(25290))))  severity failure;
	assert RAM(25291) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(25291))))  severity failure;
	assert RAM(25292) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(25292))))  severity failure;
	assert RAM(25293) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25293))))  severity failure;
	assert RAM(25294) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(25294))))  severity failure;
	assert RAM(25295) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25295))))  severity failure;
	assert RAM(25296) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(25296))))  severity failure;
	assert RAM(25297) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(25297))))  severity failure;
	assert RAM(25298) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25298))))  severity failure;
	assert RAM(25299) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25299))))  severity failure;
	assert RAM(25300) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25300))))  severity failure;
	assert RAM(25301) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(25301))))  severity failure;
	assert RAM(25302) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(25302))))  severity failure;
	assert RAM(25303) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(25303))))  severity failure;
	assert RAM(25304) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(25304))))  severity failure;
	assert RAM(25305) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(25305))))  severity failure;
	assert RAM(25306) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25306))))  severity failure;
	assert RAM(25307) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(25307))))  severity failure;
	assert RAM(25308) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25308))))  severity failure;
	assert RAM(25309) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(25309))))  severity failure;
	assert RAM(25310) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(25310))))  severity failure;
	assert RAM(25311) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25311))))  severity failure;
	assert RAM(25312) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(25312))))  severity failure;
	assert RAM(25313) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(25313))))  severity failure;
	assert RAM(25314) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(25314))))  severity failure;
	assert RAM(25315) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(25315))))  severity failure;
	assert RAM(25316) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25316))))  severity failure;
	assert RAM(25317) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(25317))))  severity failure;
	assert RAM(25318) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(25318))))  severity failure;
	assert RAM(25319) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25319))))  severity failure;
	assert RAM(25320) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25320))))  severity failure;
	assert RAM(25321) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(25321))))  severity failure;
	assert RAM(25322) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25322))))  severity failure;
	assert RAM(25323) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25323))))  severity failure;
	assert RAM(25324) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25324))))  severity failure;
	assert RAM(25325) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(25325))))  severity failure;
	assert RAM(25326) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(25326))))  severity failure;
	assert RAM(25327) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25327))))  severity failure;
	assert RAM(25328) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25328))))  severity failure;
	assert RAM(25329) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(25329))))  severity failure;
	assert RAM(25330) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25330))))  severity failure;
	assert RAM(25331) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(25331))))  severity failure;
	assert RAM(25332) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25332))))  severity failure;
	assert RAM(25333) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(25333))))  severity failure;
	assert RAM(25334) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(25334))))  severity failure;
	assert RAM(25335) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25335))))  severity failure;
	assert RAM(25336) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(25336))))  severity failure;
	assert RAM(25337) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(25337))))  severity failure;
	assert RAM(25338) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25338))))  severity failure;
	assert RAM(25339) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(25339))))  severity failure;
	assert RAM(25340) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(25340))))  severity failure;
	assert RAM(25341) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(25341))))  severity failure;
	assert RAM(25342) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(25342))))  severity failure;
	assert RAM(25343) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25343))))  severity failure;
	assert RAM(25344) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(25344))))  severity failure;
	assert RAM(25345) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(25345))))  severity failure;
	assert RAM(25346) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(25346))))  severity failure;
	assert RAM(25347) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(25347))))  severity failure;
	assert RAM(25348) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25348))))  severity failure;
	assert RAM(25349) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(25349))))  severity failure;
	assert RAM(25350) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(25350))))  severity failure;
	assert RAM(25351) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25351))))  severity failure;
	assert RAM(25352) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(25352))))  severity failure;
	assert RAM(25353) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(25353))))  severity failure;
	assert RAM(25354) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(25354))))  severity failure;
	assert RAM(25355) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25355))))  severity failure;
	assert RAM(25356) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(25356))))  severity failure;
	assert RAM(25357) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25357))))  severity failure;
	assert RAM(25358) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(25358))))  severity failure;
	assert RAM(25359) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(25359))))  severity failure;
	assert RAM(25360) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(25360))))  severity failure;
	assert RAM(25361) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(25361))))  severity failure;
	assert RAM(25362) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(25362))))  severity failure;
	assert RAM(25363) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(25363))))  severity failure;
	assert RAM(25364) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25364))))  severity failure;
	assert RAM(25365) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25365))))  severity failure;
	assert RAM(25366) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(25366))))  severity failure;
	assert RAM(25367) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(25367))))  severity failure;
	assert RAM(25368) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(25368))))  severity failure;
	assert RAM(25369) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(25369))))  severity failure;
	assert RAM(25370) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(25370))))  severity failure;
	assert RAM(25371) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25371))))  severity failure;
	assert RAM(25372) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(25372))))  severity failure;
	assert RAM(25373) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(25373))))  severity failure;
	assert RAM(25374) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(25374))))  severity failure;
	assert RAM(25375) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(25375))))  severity failure;
	assert RAM(25376) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25376))))  severity failure;
	assert RAM(25377) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25377))))  severity failure;
	assert RAM(25378) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(25378))))  severity failure;
	assert RAM(25379) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(25379))))  severity failure;
	assert RAM(25380) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25380))))  severity failure;
	assert RAM(25381) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(25381))))  severity failure;
	assert RAM(25382) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25382))))  severity failure;
	assert RAM(25383) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(25383))))  severity failure;
	assert RAM(25384) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(25384))))  severity failure;
	assert RAM(25385) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(25385))))  severity failure;
	assert RAM(25386) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(25386))))  severity failure;
	assert RAM(25387) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(25387))))  severity failure;
	assert RAM(25388) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(25388))))  severity failure;
	assert RAM(25389) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25389))))  severity failure;
	assert RAM(25390) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(25390))))  severity failure;
	assert RAM(25391) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25391))))  severity failure;
	assert RAM(25392) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25392))))  severity failure;
	assert RAM(25393) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(25393))))  severity failure;
	assert RAM(25394) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25394))))  severity failure;
	assert RAM(25395) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(25395))))  severity failure;
	assert RAM(25396) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(25396))))  severity failure;
	assert RAM(25397) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25397))))  severity failure;
	assert RAM(25398) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25398))))  severity failure;
	assert RAM(25399) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(25399))))  severity failure;
	assert RAM(25400) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25400))))  severity failure;
	assert RAM(25401) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(25401))))  severity failure;
	assert RAM(25402) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25402))))  severity failure;
	assert RAM(25403) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(25403))))  severity failure;
	assert RAM(25404) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25404))))  severity failure;
	assert RAM(25405) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(25405))))  severity failure;
	assert RAM(25406) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25406))))  severity failure;
	assert RAM(25407) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(25407))))  severity failure;
	assert RAM(25408) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(25408))))  severity failure;
	assert RAM(25409) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(25409))))  severity failure;
	assert RAM(25410) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(25410))))  severity failure;
	assert RAM(25411) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25411))))  severity failure;
	assert RAM(25412) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(25412))))  severity failure;
	assert RAM(25413) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25413))))  severity failure;
	assert RAM(25414) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(25414))))  severity failure;
	assert RAM(25415) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(25415))))  severity failure;
	assert RAM(25416) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(25416))))  severity failure;
	assert RAM(25417) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(25417))))  severity failure;
	assert RAM(25418) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(25418))))  severity failure;
	assert RAM(25419) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25419))))  severity failure;
	assert RAM(25420) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(25420))))  severity failure;
	assert RAM(25421) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(25421))))  severity failure;
	assert RAM(25422) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(25422))))  severity failure;
	assert RAM(25423) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25423))))  severity failure;
	assert RAM(25424) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(25424))))  severity failure;
	assert RAM(25425) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25425))))  severity failure;
	assert RAM(25426) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25426))))  severity failure;
	assert RAM(25427) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25427))))  severity failure;
	assert RAM(25428) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(25428))))  severity failure;
	assert RAM(25429) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(25429))))  severity failure;
	assert RAM(25430) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25430))))  severity failure;
	assert RAM(25431) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25431))))  severity failure;
	assert RAM(25432) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(25432))))  severity failure;
	assert RAM(25433) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(25433))))  severity failure;
	assert RAM(25434) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(25434))))  severity failure;
	assert RAM(25435) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25435))))  severity failure;
	assert RAM(25436) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(25436))))  severity failure;
	assert RAM(25437) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25437))))  severity failure;
	assert RAM(25438) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(25438))))  severity failure;
	assert RAM(25439) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(25439))))  severity failure;
	assert RAM(25440) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(25440))))  severity failure;
	assert RAM(25441) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25441))))  severity failure;
	assert RAM(25442) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(25442))))  severity failure;
	assert RAM(25443) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25443))))  severity failure;
	assert RAM(25444) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(25444))))  severity failure;
	assert RAM(25445) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25445))))  severity failure;
	assert RAM(25446) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(25446))))  severity failure;
	assert RAM(25447) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(25447))))  severity failure;
	assert RAM(25448) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25448))))  severity failure;
	assert RAM(25449) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(25449))))  severity failure;
	assert RAM(25450) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25450))))  severity failure;
	assert RAM(25451) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25451))))  severity failure;
	assert RAM(25452) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25452))))  severity failure;
	assert RAM(25453) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(25453))))  severity failure;
	assert RAM(25454) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(25454))))  severity failure;
	assert RAM(25455) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(25455))))  severity failure;
	assert RAM(25456) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(25456))))  severity failure;
	assert RAM(25457) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(25457))))  severity failure;
	assert RAM(25458) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(25458))))  severity failure;
	assert RAM(25459) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(25459))))  severity failure;
	assert RAM(25460) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(25460))))  severity failure;
	assert RAM(25461) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(25461))))  severity failure;
	assert RAM(25462) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(25462))))  severity failure;
	assert RAM(25463) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(25463))))  severity failure;
	assert RAM(25464) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(25464))))  severity failure;
	assert RAM(25465) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(25465))))  severity failure;
	assert RAM(25466) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25466))))  severity failure;
	assert RAM(25467) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25467))))  severity failure;
	assert RAM(25468) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25468))))  severity failure;
	assert RAM(25469) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(25469))))  severity failure;
	assert RAM(25470) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(25470))))  severity failure;
	assert RAM(25471) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(25471))))  severity failure;
	assert RAM(25472) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25472))))  severity failure;
	assert RAM(25473) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(25473))))  severity failure;
	assert RAM(25474) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(25474))))  severity failure;
	assert RAM(25475) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(25475))))  severity failure;
	assert RAM(25476) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25476))))  severity failure;
	assert RAM(25477) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(25477))))  severity failure;
	assert RAM(25478) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25478))))  severity failure;
	assert RAM(25479) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25479))))  severity failure;
	assert RAM(25480) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(25480))))  severity failure;
	assert RAM(25481) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25481))))  severity failure;
	assert RAM(25482) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(25482))))  severity failure;
	assert RAM(25483) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(25483))))  severity failure;
	assert RAM(25484) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(25484))))  severity failure;
	assert RAM(25485) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25485))))  severity failure;
	assert RAM(25486) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25486))))  severity failure;
	assert RAM(25487) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25487))))  severity failure;
	assert RAM(25488) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25488))))  severity failure;
	assert RAM(25489) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(25489))))  severity failure;
	assert RAM(25490) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(25490))))  severity failure;
	assert RAM(25491) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(25491))))  severity failure;
	assert RAM(25492) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25492))))  severity failure;
	assert RAM(25493) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(25493))))  severity failure;
	assert RAM(25494) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(25494))))  severity failure;
	assert RAM(25495) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25495))))  severity failure;
	assert RAM(25496) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25496))))  severity failure;
	assert RAM(25497) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(25497))))  severity failure;
	assert RAM(25498) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(25498))))  severity failure;
	assert RAM(25499) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(25499))))  severity failure;
	assert RAM(25500) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25500))))  severity failure;
	assert RAM(25501) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25501))))  severity failure;
	assert RAM(25502) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25502))))  severity failure;
	assert RAM(25503) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(25503))))  severity failure;
	assert RAM(25504) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25504))))  severity failure;
	assert RAM(25505) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(25505))))  severity failure;
	assert RAM(25506) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(25506))))  severity failure;
	assert RAM(25507) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(25507))))  severity failure;
	assert RAM(25508) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(25508))))  severity failure;
	assert RAM(25509) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(25509))))  severity failure;
	assert RAM(25510) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25510))))  severity failure;
	assert RAM(25511) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(25511))))  severity failure;
	assert RAM(25512) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(25512))))  severity failure;
	assert RAM(25513) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25513))))  severity failure;
	assert RAM(25514) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(25514))))  severity failure;
	assert RAM(25515) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25515))))  severity failure;
	assert RAM(25516) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(25516))))  severity failure;
	assert RAM(25517) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25517))))  severity failure;
	assert RAM(25518) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(25518))))  severity failure;
	assert RAM(25519) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(25519))))  severity failure;
	assert RAM(25520) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(25520))))  severity failure;
	assert RAM(25521) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25521))))  severity failure;
	assert RAM(25522) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25522))))  severity failure;
	assert RAM(25523) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(25523))))  severity failure;
	assert RAM(25524) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(25524))))  severity failure;
	assert RAM(25525) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25525))))  severity failure;
	assert RAM(25526) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(25526))))  severity failure;
	assert RAM(25527) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25527))))  severity failure;
	assert RAM(25528) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(25528))))  severity failure;
	assert RAM(25529) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(25529))))  severity failure;
	assert RAM(25530) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(25530))))  severity failure;
	assert RAM(25531) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25531))))  severity failure;
	assert RAM(25532) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(25532))))  severity failure;
	assert RAM(25533) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25533))))  severity failure;
	assert RAM(25534) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(25534))))  severity failure;
	assert RAM(25535) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25535))))  severity failure;
	assert RAM(25536) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25536))))  severity failure;
	assert RAM(25537) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25537))))  severity failure;
	assert RAM(25538) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(25538))))  severity failure;
	assert RAM(25539) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25539))))  severity failure;
	assert RAM(25540) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(25540))))  severity failure;
	assert RAM(25541) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25541))))  severity failure;
	assert RAM(25542) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(25542))))  severity failure;
	assert RAM(25543) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(25543))))  severity failure;
	assert RAM(25544) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(25544))))  severity failure;
	assert RAM(25545) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(25545))))  severity failure;
	assert RAM(25546) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25546))))  severity failure;
	assert RAM(25547) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25547))))  severity failure;
	assert RAM(25548) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(25548))))  severity failure;
	assert RAM(25549) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(25549))))  severity failure;
	assert RAM(25550) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25550))))  severity failure;
	assert RAM(25551) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25551))))  severity failure;
	assert RAM(25552) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25552))))  severity failure;
	assert RAM(25553) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(25553))))  severity failure;
	assert RAM(25554) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25554))))  severity failure;
	assert RAM(25555) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(25555))))  severity failure;
	assert RAM(25556) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25556))))  severity failure;
	assert RAM(25557) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25557))))  severity failure;
	assert RAM(25558) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(25558))))  severity failure;
	assert RAM(25559) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(25559))))  severity failure;
	assert RAM(25560) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25560))))  severity failure;
	assert RAM(25561) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(25561))))  severity failure;
	assert RAM(25562) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25562))))  severity failure;
	assert RAM(25563) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(25563))))  severity failure;
	assert RAM(25564) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25564))))  severity failure;
	assert RAM(25565) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(25565))))  severity failure;
	assert RAM(25566) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(25566))))  severity failure;
	assert RAM(25567) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(25567))))  severity failure;
	assert RAM(25568) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25568))))  severity failure;
	assert RAM(25569) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25569))))  severity failure;
	assert RAM(25570) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25570))))  severity failure;
	assert RAM(25571) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(25571))))  severity failure;
	assert RAM(25572) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(25572))))  severity failure;
	assert RAM(25573) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25573))))  severity failure;
	assert RAM(25574) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(25574))))  severity failure;
	assert RAM(25575) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(25575))))  severity failure;
	assert RAM(25576) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25576))))  severity failure;
	assert RAM(25577) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(25577))))  severity failure;
	assert RAM(25578) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25578))))  severity failure;
	assert RAM(25579) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(25579))))  severity failure;
	assert RAM(25580) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25580))))  severity failure;
	assert RAM(25581) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25581))))  severity failure;
	assert RAM(25582) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25582))))  severity failure;
	assert RAM(25583) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25583))))  severity failure;
	assert RAM(25584) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(25584))))  severity failure;
	assert RAM(25585) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(25585))))  severity failure;
	assert RAM(25586) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(25586))))  severity failure;
	assert RAM(25587) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(25587))))  severity failure;
	assert RAM(25588) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(25588))))  severity failure;
	assert RAM(25589) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(25589))))  severity failure;
	assert RAM(25590) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(25590))))  severity failure;
	assert RAM(25591) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(25591))))  severity failure;
	assert RAM(25592) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(25592))))  severity failure;
	assert RAM(25593) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(25593))))  severity failure;
	assert RAM(25594) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(25594))))  severity failure;
	assert RAM(25595) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25595))))  severity failure;
	assert RAM(25596) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25596))))  severity failure;
	assert RAM(25597) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25597))))  severity failure;
	assert RAM(25598) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(25598))))  severity failure;
	assert RAM(25599) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(25599))))  severity failure;
	assert RAM(25600) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(25600))))  severity failure;
	assert RAM(25601) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(25601))))  severity failure;
	assert RAM(25602) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(25602))))  severity failure;
	assert RAM(25603) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(25603))))  severity failure;
	assert RAM(25604) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25604))))  severity failure;
	assert RAM(25605) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(25605))))  severity failure;
	assert RAM(25606) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(25606))))  severity failure;
	assert RAM(25607) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(25607))))  severity failure;
	assert RAM(25608) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(25608))))  severity failure;
	assert RAM(25609) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(25609))))  severity failure;
	assert RAM(25610) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25610))))  severity failure;
	assert RAM(25611) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(25611))))  severity failure;
	assert RAM(25612) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(25612))))  severity failure;
	assert RAM(25613) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25613))))  severity failure;
	assert RAM(25614) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25614))))  severity failure;
	assert RAM(25615) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25615))))  severity failure;
	assert RAM(25616) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25616))))  severity failure;
	assert RAM(25617) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25617))))  severity failure;
	assert RAM(25618) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(25618))))  severity failure;
	assert RAM(25619) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(25619))))  severity failure;
	assert RAM(25620) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(25620))))  severity failure;
	assert RAM(25621) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25621))))  severity failure;
	assert RAM(25622) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25622))))  severity failure;
	assert RAM(25623) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(25623))))  severity failure;
	assert RAM(25624) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(25624))))  severity failure;
	assert RAM(25625) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(25625))))  severity failure;
	assert RAM(25626) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(25626))))  severity failure;
	assert RAM(25627) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(25627))))  severity failure;
	assert RAM(25628) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(25628))))  severity failure;
	assert RAM(25629) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(25629))))  severity failure;
	assert RAM(25630) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(25630))))  severity failure;
	assert RAM(25631) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(25631))))  severity failure;
	assert RAM(25632) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(25632))))  severity failure;
	assert RAM(25633) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(25633))))  severity failure;
	assert RAM(25634) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25634))))  severity failure;
	assert RAM(25635) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(25635))))  severity failure;
	assert RAM(25636) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(25636))))  severity failure;
	assert RAM(25637) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(25637))))  severity failure;
	assert RAM(25638) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(25638))))  severity failure;
	assert RAM(25639) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(25639))))  severity failure;
	assert RAM(25640) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(25640))))  severity failure;
	assert RAM(25641) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(25641))))  severity failure;
	assert RAM(25642) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(25642))))  severity failure;
	assert RAM(25643) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(25643))))  severity failure;
	assert RAM(25644) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(25644))))  severity failure;
	assert RAM(25645) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25645))))  severity failure;
	assert RAM(25646) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(25646))))  severity failure;
	assert RAM(25647) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25647))))  severity failure;
	assert RAM(25648) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(25648))))  severity failure;
	assert RAM(25649) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(25649))))  severity failure;
	assert RAM(25650) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(25650))))  severity failure;
	assert RAM(25651) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25651))))  severity failure;
	assert RAM(25652) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(25652))))  severity failure;
	assert RAM(25653) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25653))))  severity failure;
	assert RAM(25654) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(25654))))  severity failure;
	assert RAM(25655) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25655))))  severity failure;
	assert RAM(25656) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(25656))))  severity failure;
	assert RAM(25657) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(25657))))  severity failure;
	assert RAM(25658) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(25658))))  severity failure;
	assert RAM(25659) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(25659))))  severity failure;
	assert RAM(25660) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(25660))))  severity failure;
	assert RAM(25661) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25661))))  severity failure;
	assert RAM(25662) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(25662))))  severity failure;
	assert RAM(25663) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(25663))))  severity failure;
	assert RAM(25664) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25664))))  severity failure;
	assert RAM(25665) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(25665))))  severity failure;
	assert RAM(25666) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(25666))))  severity failure;
	assert RAM(25667) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(25667))))  severity failure;
	assert RAM(25668) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25668))))  severity failure;
	assert RAM(25669) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25669))))  severity failure;
	assert RAM(25670) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(25670))))  severity failure;
	assert RAM(25671) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(25671))))  severity failure;
	assert RAM(25672) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25672))))  severity failure;
	assert RAM(25673) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25673))))  severity failure;
	assert RAM(25674) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(25674))))  severity failure;
	assert RAM(25675) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(25675))))  severity failure;
	assert RAM(25676) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25676))))  severity failure;
	assert RAM(25677) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25677))))  severity failure;
	assert RAM(25678) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(25678))))  severity failure;
	assert RAM(25679) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(25679))))  severity failure;
	assert RAM(25680) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(25680))))  severity failure;
	assert RAM(25681) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(25681))))  severity failure;
	assert RAM(25682) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(25682))))  severity failure;
	assert RAM(25683) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25683))))  severity failure;
	assert RAM(25684) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(25684))))  severity failure;
	assert RAM(25685) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25685))))  severity failure;
	assert RAM(25686) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(25686))))  severity failure;
	assert RAM(25687) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(25687))))  severity failure;
	assert RAM(25688) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(25688))))  severity failure;
	assert RAM(25689) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(25689))))  severity failure;
	assert RAM(25690) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(25690))))  severity failure;
	assert RAM(25691) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25691))))  severity failure;
	assert RAM(25692) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25692))))  severity failure;
	assert RAM(25693) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(25693))))  severity failure;
	assert RAM(25694) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(25694))))  severity failure;
	assert RAM(25695) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25695))))  severity failure;
	assert RAM(25696) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(25696))))  severity failure;
	assert RAM(25697) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25697))))  severity failure;
	assert RAM(25698) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(25698))))  severity failure;
	assert RAM(25699) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25699))))  severity failure;
	assert RAM(25700) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(25700))))  severity failure;
	assert RAM(25701) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(25701))))  severity failure;
	assert RAM(25702) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(25702))))  severity failure;
	assert RAM(25703) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(25703))))  severity failure;
	assert RAM(25704) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(25704))))  severity failure;
	assert RAM(25705) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(25705))))  severity failure;
	assert RAM(25706) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(25706))))  severity failure;
	assert RAM(25707) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(25707))))  severity failure;
	assert RAM(25708) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(25708))))  severity failure;
	assert RAM(25709) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(25709))))  severity failure;
	assert RAM(25710) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(25710))))  severity failure;
	assert RAM(25711) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(25711))))  severity failure;
	assert RAM(25712) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25712))))  severity failure;
	assert RAM(25713) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(25713))))  severity failure;
	assert RAM(25714) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25714))))  severity failure;
	assert RAM(25715) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(25715))))  severity failure;
	assert RAM(25716) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(25716))))  severity failure;
	assert RAM(25717) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25717))))  severity failure;
	assert RAM(25718) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25718))))  severity failure;
	assert RAM(25719) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25719))))  severity failure;
	assert RAM(25720) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(25720))))  severity failure;
	assert RAM(25721) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(25721))))  severity failure;
	assert RAM(25722) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(25722))))  severity failure;
	assert RAM(25723) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(25723))))  severity failure;
	assert RAM(25724) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(25724))))  severity failure;
	assert RAM(25725) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(25725))))  severity failure;
	assert RAM(25726) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25726))))  severity failure;
	assert RAM(25727) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25727))))  severity failure;
	assert RAM(25728) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(25728))))  severity failure;
	assert RAM(25729) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(25729))))  severity failure;
	assert RAM(25730) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(25730))))  severity failure;
	assert RAM(25731) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(25731))))  severity failure;
	assert RAM(25732) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(25732))))  severity failure;
	assert RAM(25733) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(25733))))  severity failure;
	assert RAM(25734) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(25734))))  severity failure;
	assert RAM(25735) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25735))))  severity failure;
	assert RAM(25736) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25736))))  severity failure;
	assert RAM(25737) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25737))))  severity failure;
	assert RAM(25738) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25738))))  severity failure;
	assert RAM(25739) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(25739))))  severity failure;
	assert RAM(25740) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25740))))  severity failure;
	assert RAM(25741) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(25741))))  severity failure;
	assert RAM(25742) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(25742))))  severity failure;
	assert RAM(25743) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25743))))  severity failure;
	assert RAM(25744) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25744))))  severity failure;
	assert RAM(25745) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(25745))))  severity failure;
	assert RAM(25746) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25746))))  severity failure;
	assert RAM(25747) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(25747))))  severity failure;
	assert RAM(25748) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(25748))))  severity failure;
	assert RAM(25749) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25749))))  severity failure;
	assert RAM(25750) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(25750))))  severity failure;
	assert RAM(25751) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25751))))  severity failure;
	assert RAM(25752) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(25752))))  severity failure;
	assert RAM(25753) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(25753))))  severity failure;
	assert RAM(25754) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(25754))))  severity failure;
	assert RAM(25755) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(25755))))  severity failure;
	assert RAM(25756) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(25756))))  severity failure;
	assert RAM(25757) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25757))))  severity failure;
	assert RAM(25758) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(25758))))  severity failure;
	assert RAM(25759) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(25759))))  severity failure;
	assert RAM(25760) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(25760))))  severity failure;
	assert RAM(25761) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(25761))))  severity failure;
	assert RAM(25762) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(25762))))  severity failure;
	assert RAM(25763) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(25763))))  severity failure;
	assert RAM(25764) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25764))))  severity failure;
	assert RAM(25765) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(25765))))  severity failure;
	assert RAM(25766) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(25766))))  severity failure;
	assert RAM(25767) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(25767))))  severity failure;
	assert RAM(25768) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(25768))))  severity failure;
	assert RAM(25769) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(25769))))  severity failure;
	assert RAM(25770) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(25770))))  severity failure;
	assert RAM(25771) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25771))))  severity failure;
	assert RAM(25772) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(25772))))  severity failure;
	assert RAM(25773) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(25773))))  severity failure;
	assert RAM(25774) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25774))))  severity failure;
	assert RAM(25775) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(25775))))  severity failure;
	assert RAM(25776) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(25776))))  severity failure;
	assert RAM(25777) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(25777))))  severity failure;
	assert RAM(25778) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25778))))  severity failure;
	assert RAM(25779) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25779))))  severity failure;
	assert RAM(25780) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25780))))  severity failure;
	assert RAM(25781) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(25781))))  severity failure;
	assert RAM(25782) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25782))))  severity failure;
	assert RAM(25783) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25783))))  severity failure;
	assert RAM(25784) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25784))))  severity failure;
	assert RAM(25785) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(25785))))  severity failure;
	assert RAM(25786) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(25786))))  severity failure;
	assert RAM(25787) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25787))))  severity failure;
	assert RAM(25788) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25788))))  severity failure;
	assert RAM(25789) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(25789))))  severity failure;
	assert RAM(25790) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(25790))))  severity failure;
	assert RAM(25791) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(25791))))  severity failure;
	assert RAM(25792) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25792))))  severity failure;
	assert RAM(25793) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(25793))))  severity failure;
	assert RAM(25794) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(25794))))  severity failure;
	assert RAM(25795) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(25795))))  severity failure;
	assert RAM(25796) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25796))))  severity failure;
	assert RAM(25797) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(25797))))  severity failure;
	assert RAM(25798) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25798))))  severity failure;
	assert RAM(25799) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(25799))))  severity failure;
	assert RAM(25800) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(25800))))  severity failure;
	assert RAM(25801) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(25801))))  severity failure;
	assert RAM(25802) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(25802))))  severity failure;
	assert RAM(25803) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(25803))))  severity failure;
	assert RAM(25804) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25804))))  severity failure;
	assert RAM(25805) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(25805))))  severity failure;
	assert RAM(25806) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(25806))))  severity failure;
	assert RAM(25807) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(25807))))  severity failure;
	assert RAM(25808) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25808))))  severity failure;
	assert RAM(25809) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(25809))))  severity failure;
	assert RAM(25810) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(25810))))  severity failure;
	assert RAM(25811) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(25811))))  severity failure;
	assert RAM(25812) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(25812))))  severity failure;
	assert RAM(25813) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(25813))))  severity failure;
	assert RAM(25814) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(25814))))  severity failure;
	assert RAM(25815) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(25815))))  severity failure;
	assert RAM(25816) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25816))))  severity failure;
	assert RAM(25817) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25817))))  severity failure;
	assert RAM(25818) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(25818))))  severity failure;
	assert RAM(25819) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25819))))  severity failure;
	assert RAM(25820) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(25820))))  severity failure;
	assert RAM(25821) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(25821))))  severity failure;
	assert RAM(25822) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(25822))))  severity failure;
	assert RAM(25823) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(25823))))  severity failure;
	assert RAM(25824) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25824))))  severity failure;
	assert RAM(25825) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(25825))))  severity failure;
	assert RAM(25826) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(25826))))  severity failure;
	assert RAM(25827) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(25827))))  severity failure;
	assert RAM(25828) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(25828))))  severity failure;
	assert RAM(25829) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(25829))))  severity failure;
	assert RAM(25830) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25830))))  severity failure;
	assert RAM(25831) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(25831))))  severity failure;
	assert RAM(25832) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(25832))))  severity failure;
	assert RAM(25833) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(25833))))  severity failure;
	assert RAM(25834) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(25834))))  severity failure;
	assert RAM(25835) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(25835))))  severity failure;
	assert RAM(25836) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(25836))))  severity failure;
	assert RAM(25837) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(25837))))  severity failure;
	assert RAM(25838) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(25838))))  severity failure;
	assert RAM(25839) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(25839))))  severity failure;
	assert RAM(25840) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25840))))  severity failure;
	assert RAM(25841) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(25841))))  severity failure;
	assert RAM(25842) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25842))))  severity failure;
	assert RAM(25843) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25843))))  severity failure;
	assert RAM(25844) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(25844))))  severity failure;
	assert RAM(25845) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(25845))))  severity failure;
	assert RAM(25846) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(25846))))  severity failure;
	assert RAM(25847) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(25847))))  severity failure;
	assert RAM(25848) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(25848))))  severity failure;
	assert RAM(25849) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(25849))))  severity failure;
	assert RAM(25850) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25850))))  severity failure;
	assert RAM(25851) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25851))))  severity failure;
	assert RAM(25852) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(25852))))  severity failure;
	assert RAM(25853) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(25853))))  severity failure;
	assert RAM(25854) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(25854))))  severity failure;
	assert RAM(25855) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(25855))))  severity failure;
	assert RAM(25856) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(25856))))  severity failure;
	assert RAM(25857) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(25857))))  severity failure;
	assert RAM(25858) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(25858))))  severity failure;
	assert RAM(25859) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(25859))))  severity failure;
	assert RAM(25860) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25860))))  severity failure;
	assert RAM(25861) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25861))))  severity failure;
	assert RAM(25862) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(25862))))  severity failure;
	assert RAM(25863) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(25863))))  severity failure;
	assert RAM(25864) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(25864))))  severity failure;
	assert RAM(25865) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(25865))))  severity failure;
	assert RAM(25866) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(25866))))  severity failure;
	assert RAM(25867) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(25867))))  severity failure;
	assert RAM(25868) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(25868))))  severity failure;
	assert RAM(25869) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(25869))))  severity failure;
	assert RAM(25870) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(25870))))  severity failure;
	assert RAM(25871) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(25871))))  severity failure;
	assert RAM(25872) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(25872))))  severity failure;
	assert RAM(25873) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(25873))))  severity failure;
	assert RAM(25874) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(25874))))  severity failure;
	assert RAM(25875) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(25875))))  severity failure;
	assert RAM(25876) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(25876))))  severity failure;
	assert RAM(25877) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(25877))))  severity failure;
	assert RAM(25878) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(25878))))  severity failure;
	assert RAM(25879) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(25879))))  severity failure;
	assert RAM(25880) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(25880))))  severity failure;
	assert RAM(25881) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(25881))))  severity failure;
	assert RAM(25882) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(25882))))  severity failure;
	assert RAM(25883) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25883))))  severity failure;
	assert RAM(25884) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(25884))))  severity failure;
	assert RAM(25885) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(25885))))  severity failure;
	assert RAM(25886) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(25886))))  severity failure;
	assert RAM(25887) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(25887))))  severity failure;
	assert RAM(25888) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(25888))))  severity failure;
	assert RAM(25889) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25889))))  severity failure;
	assert RAM(25890) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(25890))))  severity failure;
	assert RAM(25891) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25891))))  severity failure;
	assert RAM(25892) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(25892))))  severity failure;
	assert RAM(25893) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(25893))))  severity failure;
	assert RAM(25894) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(25894))))  severity failure;
	assert RAM(25895) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(25895))))  severity failure;
	assert RAM(25896) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25896))))  severity failure;
	assert RAM(25897) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(25897))))  severity failure;
	assert RAM(25898) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(25898))))  severity failure;
	assert RAM(25899) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(25899))))  severity failure;
	assert RAM(25900) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(25900))))  severity failure;
	assert RAM(25901) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25901))))  severity failure;
	assert RAM(25902) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(25902))))  severity failure;
	assert RAM(25903) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(25903))))  severity failure;
	assert RAM(25904) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(25904))))  severity failure;
	assert RAM(25905) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25905))))  severity failure;
	assert RAM(25906) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(25906))))  severity failure;
	assert RAM(25907) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(25907))))  severity failure;
	assert RAM(25908) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(25908))))  severity failure;
	assert RAM(25909) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(25909))))  severity failure;
	assert RAM(25910) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(25910))))  severity failure;
	assert RAM(25911) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(25911))))  severity failure;
	assert RAM(25912) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(25912))))  severity failure;
	assert RAM(25913) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(25913))))  severity failure;
	assert RAM(25914) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25914))))  severity failure;
	assert RAM(25915) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(25915))))  severity failure;
	assert RAM(25916) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(25916))))  severity failure;
	assert RAM(25917) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(25917))))  severity failure;
	assert RAM(25918) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(25918))))  severity failure;
	assert RAM(25919) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(25919))))  severity failure;
	assert RAM(25920) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(25920))))  severity failure;
	assert RAM(25921) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(25921))))  severity failure;
	assert RAM(25922) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(25922))))  severity failure;
	assert RAM(25923) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(25923))))  severity failure;
	assert RAM(25924) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(25924))))  severity failure;
	assert RAM(25925) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(25925))))  severity failure;
	assert RAM(25926) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(25926))))  severity failure;
	assert RAM(25927) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(25927))))  severity failure;
	assert RAM(25928) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(25928))))  severity failure;
	assert RAM(25929) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(25929))))  severity failure;
	assert RAM(25930) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(25930))))  severity failure;
	assert RAM(25931) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(25931))))  severity failure;
	assert RAM(25932) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25932))))  severity failure;
	assert RAM(25933) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(25933))))  severity failure;
	assert RAM(25934) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(25934))))  severity failure;
	assert RAM(25935) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(25935))))  severity failure;
	assert RAM(25936) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(25936))))  severity failure;
	assert RAM(25937) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(25937))))  severity failure;
	assert RAM(25938) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(25938))))  severity failure;
	assert RAM(25939) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(25939))))  severity failure;
	assert RAM(25940) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(25940))))  severity failure;
	assert RAM(25941) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(25941))))  severity failure;
	assert RAM(25942) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(25942))))  severity failure;
	assert RAM(25943) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(25943))))  severity failure;
	assert RAM(25944) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(25944))))  severity failure;
	assert RAM(25945) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(25945))))  severity failure;
	assert RAM(25946) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(25946))))  severity failure;
	assert RAM(25947) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(25947))))  severity failure;
	assert RAM(25948) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(25948))))  severity failure;
	assert RAM(25949) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(25949))))  severity failure;
	assert RAM(25950) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(25950))))  severity failure;
	assert RAM(25951) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25951))))  severity failure;
	assert RAM(25952) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(25952))))  severity failure;
	assert RAM(25953) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(25953))))  severity failure;
	assert RAM(25954) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(25954))))  severity failure;
	assert RAM(25955) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(25955))))  severity failure;
	assert RAM(25956) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25956))))  severity failure;
	assert RAM(25957) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(25957))))  severity failure;
	assert RAM(25958) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(25958))))  severity failure;
	assert RAM(25959) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(25959))))  severity failure;
	assert RAM(25960) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(25960))))  severity failure;
	assert RAM(25961) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(25961))))  severity failure;
	assert RAM(25962) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(25962))))  severity failure;
	assert RAM(25963) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(25963))))  severity failure;
	assert RAM(25964) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(25964))))  severity failure;
	assert RAM(25965) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(25965))))  severity failure;
	assert RAM(25966) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(25966))))  severity failure;
	assert RAM(25967) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(25967))))  severity failure;
	assert RAM(25968) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(25968))))  severity failure;
	assert RAM(25969) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(25969))))  severity failure;
	assert RAM(25970) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(25970))))  severity failure;
	assert RAM(25971) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(25971))))  severity failure;
	assert RAM(25972) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(25972))))  severity failure;
	assert RAM(25973) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(25973))))  severity failure;
	assert RAM(25974) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(25974))))  severity failure;
	assert RAM(25975) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(25975))))  severity failure;
	assert RAM(25976) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(25976))))  severity failure;
	assert RAM(25977) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(25977))))  severity failure;
	assert RAM(25978) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(25978))))  severity failure;
	assert RAM(25979) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(25979))))  severity failure;
	assert RAM(25980) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(25980))))  severity failure;
	assert RAM(25981) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(25981))))  severity failure;
	assert RAM(25982) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(25982))))  severity failure;
	assert RAM(25983) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(25983))))  severity failure;
	assert RAM(25984) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(25984))))  severity failure;
	assert RAM(25985) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(25985))))  severity failure;
	assert RAM(25986) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(25986))))  severity failure;
	assert RAM(25987) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(25987))))  severity failure;
	assert RAM(25988) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(25988))))  severity failure;
	assert RAM(25989) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(25989))))  severity failure;
	assert RAM(25990) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(25990))))  severity failure;
	assert RAM(25991) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(25991))))  severity failure;
	assert RAM(25992) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(25992))))  severity failure;
	assert RAM(25993) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(25993))))  severity failure;
	assert RAM(25994) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(25994))))  severity failure;
	assert RAM(25995) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(25995))))  severity failure;
	assert RAM(25996) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(25996))))  severity failure;
	assert RAM(25997) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(25997))))  severity failure;
	assert RAM(25998) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(25998))))  severity failure;
	assert RAM(25999) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(25999))))  severity failure;
	assert RAM(26000) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(26000))))  severity failure;
	assert RAM(26001) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(26001))))  severity failure;
	assert RAM(26002) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(26002))))  severity failure;
	assert RAM(26003) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(26003))))  severity failure;
	assert RAM(26004) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(26004))))  severity failure;
	assert RAM(26005) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(26005))))  severity failure;
	assert RAM(26006) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26006))))  severity failure;
	assert RAM(26007) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26007))))  severity failure;
	assert RAM(26008) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26008))))  severity failure;
	assert RAM(26009) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(26009))))  severity failure;
	assert RAM(26010) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(26010))))  severity failure;
	assert RAM(26011) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(26011))))  severity failure;
	assert RAM(26012) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(26012))))  severity failure;
	assert RAM(26013) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(26013))))  severity failure;
	assert RAM(26014) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26014))))  severity failure;
	assert RAM(26015) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(26015))))  severity failure;
	assert RAM(26016) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(26016))))  severity failure;
	assert RAM(26017) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(26017))))  severity failure;
	assert RAM(26018) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(26018))))  severity failure;
	assert RAM(26019) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26019))))  severity failure;
	assert RAM(26020) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(26020))))  severity failure;
	assert RAM(26021) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(26021))))  severity failure;
	assert RAM(26022) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26022))))  severity failure;
	assert RAM(26023) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(26023))))  severity failure;
	assert RAM(26024) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26024))))  severity failure;
	assert RAM(26025) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(26025))))  severity failure;
	assert RAM(26026) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(26026))))  severity failure;
	assert RAM(26027) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(26027))))  severity failure;
	assert RAM(26028) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(26028))))  severity failure;
	assert RAM(26029) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(26029))))  severity failure;
	assert RAM(26030) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26030))))  severity failure;
	assert RAM(26031) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(26031))))  severity failure;
	assert RAM(26032) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26032))))  severity failure;
	assert RAM(26033) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(26033))))  severity failure;
	assert RAM(26034) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(26034))))  severity failure;
	assert RAM(26035) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26035))))  severity failure;
	assert RAM(26036) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(26036))))  severity failure;
	assert RAM(26037) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(26037))))  severity failure;
	assert RAM(26038) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26038))))  severity failure;
	assert RAM(26039) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(26039))))  severity failure;
	assert RAM(26040) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(26040))))  severity failure;
	assert RAM(26041) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26041))))  severity failure;
	assert RAM(26042) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26042))))  severity failure;
	assert RAM(26043) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(26043))))  severity failure;
	assert RAM(26044) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26044))))  severity failure;
	assert RAM(26045) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26045))))  severity failure;
	assert RAM(26046) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26046))))  severity failure;
	assert RAM(26047) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26047))))  severity failure;
	assert RAM(26048) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(26048))))  severity failure;
	assert RAM(26049) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(26049))))  severity failure;
	assert RAM(26050) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(26050))))  severity failure;
	assert RAM(26051) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(26051))))  severity failure;
	assert RAM(26052) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(26052))))  severity failure;
	assert RAM(26053) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(26053))))  severity failure;
	assert RAM(26054) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26054))))  severity failure;
	assert RAM(26055) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(26055))))  severity failure;
	assert RAM(26056) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(26056))))  severity failure;
	assert RAM(26057) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(26057))))  severity failure;
	assert RAM(26058) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(26058))))  severity failure;
	assert RAM(26059) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26059))))  severity failure;
	assert RAM(26060) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26060))))  severity failure;
	assert RAM(26061) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26061))))  severity failure;
	assert RAM(26062) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(26062))))  severity failure;
	assert RAM(26063) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(26063))))  severity failure;
	assert RAM(26064) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(26064))))  severity failure;
	assert RAM(26065) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(26065))))  severity failure;
	assert RAM(26066) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(26066))))  severity failure;
	assert RAM(26067) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(26067))))  severity failure;
	assert RAM(26068) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(26068))))  severity failure;
	assert RAM(26069) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(26069))))  severity failure;
	assert RAM(26070) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26070))))  severity failure;
	assert RAM(26071) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(26071))))  severity failure;
	assert RAM(26072) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(26072))))  severity failure;
	assert RAM(26073) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26073))))  severity failure;
	assert RAM(26074) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(26074))))  severity failure;
	assert RAM(26075) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26075))))  severity failure;
	assert RAM(26076) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(26076))))  severity failure;
	assert RAM(26077) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(26077))))  severity failure;
	assert RAM(26078) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(26078))))  severity failure;
	assert RAM(26079) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(26079))))  severity failure;
	assert RAM(26080) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26080))))  severity failure;
	assert RAM(26081) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(26081))))  severity failure;
	assert RAM(26082) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26082))))  severity failure;
	assert RAM(26083) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(26083))))  severity failure;
	assert RAM(26084) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(26084))))  severity failure;
	assert RAM(26085) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(26085))))  severity failure;
	assert RAM(26086) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(26086))))  severity failure;
	assert RAM(26087) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26087))))  severity failure;
	assert RAM(26088) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(26088))))  severity failure;
	assert RAM(26089) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(26089))))  severity failure;
	assert RAM(26090) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26090))))  severity failure;
	assert RAM(26091) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26091))))  severity failure;
	assert RAM(26092) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(26092))))  severity failure;
	assert RAM(26093) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26093))))  severity failure;
	assert RAM(26094) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(26094))))  severity failure;
	assert RAM(26095) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(26095))))  severity failure;
	assert RAM(26096) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26096))))  severity failure;
	assert RAM(26097) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(26097))))  severity failure;
	assert RAM(26098) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(26098))))  severity failure;
	assert RAM(26099) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26099))))  severity failure;
	assert RAM(26100) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(26100))))  severity failure;
	assert RAM(26101) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26101))))  severity failure;
	assert RAM(26102) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(26102))))  severity failure;
	assert RAM(26103) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(26103))))  severity failure;
	assert RAM(26104) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(26104))))  severity failure;
	assert RAM(26105) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(26105))))  severity failure;
	assert RAM(26106) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(26106))))  severity failure;
	assert RAM(26107) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26107))))  severity failure;
	assert RAM(26108) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(26108))))  severity failure;
	assert RAM(26109) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(26109))))  severity failure;
	assert RAM(26110) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26110))))  severity failure;
	assert RAM(26111) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26111))))  severity failure;
	assert RAM(26112) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(26112))))  severity failure;
	assert RAM(26113) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26113))))  severity failure;
	assert RAM(26114) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26114))))  severity failure;
	assert RAM(26115) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(26115))))  severity failure;
	assert RAM(26116) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26116))))  severity failure;
	assert RAM(26117) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26117))))  severity failure;
	assert RAM(26118) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26118))))  severity failure;
	assert RAM(26119) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(26119))))  severity failure;
	assert RAM(26120) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26120))))  severity failure;
	assert RAM(26121) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(26121))))  severity failure;
	assert RAM(26122) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(26122))))  severity failure;
	assert RAM(26123) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(26123))))  severity failure;
	assert RAM(26124) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(26124))))  severity failure;
	assert RAM(26125) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26125))))  severity failure;
	assert RAM(26126) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(26126))))  severity failure;
	assert RAM(26127) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(26127))))  severity failure;
	assert RAM(26128) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26128))))  severity failure;
	assert RAM(26129) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(26129))))  severity failure;
	assert RAM(26130) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(26130))))  severity failure;
	assert RAM(26131) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(26131))))  severity failure;
	assert RAM(26132) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26132))))  severity failure;
	assert RAM(26133) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(26133))))  severity failure;
	assert RAM(26134) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(26134))))  severity failure;
	assert RAM(26135) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(26135))))  severity failure;
	assert RAM(26136) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(26136))))  severity failure;
	assert RAM(26137) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26137))))  severity failure;
	assert RAM(26138) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(26138))))  severity failure;
	assert RAM(26139) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(26139))))  severity failure;
	assert RAM(26140) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(26140))))  severity failure;
	assert RAM(26141) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(26141))))  severity failure;
	assert RAM(26142) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(26142))))  severity failure;
	assert RAM(26143) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(26143))))  severity failure;
	assert RAM(26144) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26144))))  severity failure;
	assert RAM(26145) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26145))))  severity failure;
	assert RAM(26146) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(26146))))  severity failure;
	assert RAM(26147) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(26147))))  severity failure;
	assert RAM(26148) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(26148))))  severity failure;
	assert RAM(26149) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26149))))  severity failure;
	assert RAM(26150) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(26150))))  severity failure;
	assert RAM(26151) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26151))))  severity failure;
	assert RAM(26152) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26152))))  severity failure;
	assert RAM(26153) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26153))))  severity failure;
	assert RAM(26154) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(26154))))  severity failure;
	assert RAM(26155) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26155))))  severity failure;
	assert RAM(26156) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26156))))  severity failure;
	assert RAM(26157) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(26157))))  severity failure;
	assert RAM(26158) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26158))))  severity failure;
	assert RAM(26159) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(26159))))  severity failure;
	assert RAM(26160) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(26160))))  severity failure;
	assert RAM(26161) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26161))))  severity failure;
	assert RAM(26162) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26162))))  severity failure;
	assert RAM(26163) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(26163))))  severity failure;
	assert RAM(26164) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(26164))))  severity failure;
	assert RAM(26165) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26165))))  severity failure;
	assert RAM(26166) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(26166))))  severity failure;
	assert RAM(26167) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(26167))))  severity failure;
	assert RAM(26168) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(26168))))  severity failure;
	assert RAM(26169) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(26169))))  severity failure;
	assert RAM(26170) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(26170))))  severity failure;
	assert RAM(26171) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(26171))))  severity failure;
	assert RAM(26172) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(26172))))  severity failure;
	assert RAM(26173) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(26173))))  severity failure;
	assert RAM(26174) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26174))))  severity failure;
	assert RAM(26175) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(26175))))  severity failure;
	assert RAM(26176) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(26176))))  severity failure;
	assert RAM(26177) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(26177))))  severity failure;
	assert RAM(26178) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26178))))  severity failure;
	assert RAM(26179) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(26179))))  severity failure;
	assert RAM(26180) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(26180))))  severity failure;
	assert RAM(26181) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26181))))  severity failure;
	assert RAM(26182) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(26182))))  severity failure;
	assert RAM(26183) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(26183))))  severity failure;
	assert RAM(26184) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(26184))))  severity failure;
	assert RAM(26185) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26185))))  severity failure;
	assert RAM(26186) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(26186))))  severity failure;
	assert RAM(26187) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(26187))))  severity failure;
	assert RAM(26188) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(26188))))  severity failure;
	assert RAM(26189) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26189))))  severity failure;
	assert RAM(26190) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(26190))))  severity failure;
	assert RAM(26191) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(26191))))  severity failure;
	assert RAM(26192) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(26192))))  severity failure;
	assert RAM(26193) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(26193))))  severity failure;
	assert RAM(26194) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26194))))  severity failure;
	assert RAM(26195) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26195))))  severity failure;
	assert RAM(26196) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(26196))))  severity failure;
	assert RAM(26197) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26197))))  severity failure;
	assert RAM(26198) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26198))))  severity failure;
	assert RAM(26199) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(26199))))  severity failure;
	assert RAM(26200) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(26200))))  severity failure;
	assert RAM(26201) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26201))))  severity failure;
	assert RAM(26202) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(26202))))  severity failure;
	assert RAM(26203) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26203))))  severity failure;
	assert RAM(26204) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26204))))  severity failure;
	assert RAM(26205) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26205))))  severity failure;
	assert RAM(26206) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26206))))  severity failure;
	assert RAM(26207) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(26207))))  severity failure;
	assert RAM(26208) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26208))))  severity failure;
	assert RAM(26209) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(26209))))  severity failure;
	assert RAM(26210) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(26210))))  severity failure;
	assert RAM(26211) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(26211))))  severity failure;
	assert RAM(26212) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(26212))))  severity failure;
	assert RAM(26213) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(26213))))  severity failure;
	assert RAM(26214) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(26214))))  severity failure;
	assert RAM(26215) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26215))))  severity failure;
	assert RAM(26216) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(26216))))  severity failure;
	assert RAM(26217) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26217))))  severity failure;
	assert RAM(26218) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(26218))))  severity failure;
	assert RAM(26219) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(26219))))  severity failure;
	assert RAM(26220) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26220))))  severity failure;
	assert RAM(26221) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(26221))))  severity failure;
	assert RAM(26222) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(26222))))  severity failure;
	assert RAM(26223) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(26223))))  severity failure;
	assert RAM(26224) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(26224))))  severity failure;
	assert RAM(26225) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26225))))  severity failure;
	assert RAM(26226) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(26226))))  severity failure;
	assert RAM(26227) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26227))))  severity failure;
	assert RAM(26228) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26228))))  severity failure;
	assert RAM(26229) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26229))))  severity failure;
	assert RAM(26230) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26230))))  severity failure;
	assert RAM(26231) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(26231))))  severity failure;
	assert RAM(26232) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(26232))))  severity failure;
	assert RAM(26233) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(26233))))  severity failure;
	assert RAM(26234) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26234))))  severity failure;
	assert RAM(26235) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(26235))))  severity failure;
	assert RAM(26236) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(26236))))  severity failure;
	assert RAM(26237) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(26237))))  severity failure;
	assert RAM(26238) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(26238))))  severity failure;
	assert RAM(26239) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(26239))))  severity failure;
	assert RAM(26240) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(26240))))  severity failure;
	assert RAM(26241) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(26241))))  severity failure;
	assert RAM(26242) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(26242))))  severity failure;
	assert RAM(26243) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(26243))))  severity failure;
	assert RAM(26244) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(26244))))  severity failure;
	assert RAM(26245) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26245))))  severity failure;
	assert RAM(26246) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26246))))  severity failure;
	assert RAM(26247) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(26247))))  severity failure;
	assert RAM(26248) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(26248))))  severity failure;
	assert RAM(26249) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(26249))))  severity failure;
	assert RAM(26250) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26250))))  severity failure;
	assert RAM(26251) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(26251))))  severity failure;
	assert RAM(26252) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(26252))))  severity failure;
	assert RAM(26253) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(26253))))  severity failure;
	assert RAM(26254) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26254))))  severity failure;
	assert RAM(26255) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(26255))))  severity failure;
	assert RAM(26256) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(26256))))  severity failure;
	assert RAM(26257) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(26257))))  severity failure;
	assert RAM(26258) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(26258))))  severity failure;
	assert RAM(26259) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26259))))  severity failure;
	assert RAM(26260) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(26260))))  severity failure;
	assert RAM(26261) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26261))))  severity failure;
	assert RAM(26262) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(26262))))  severity failure;
	assert RAM(26263) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26263))))  severity failure;
	assert RAM(26264) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(26264))))  severity failure;
	assert RAM(26265) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(26265))))  severity failure;
	assert RAM(26266) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(26266))))  severity failure;
	assert RAM(26267) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26267))))  severity failure;
	assert RAM(26268) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(26268))))  severity failure;
	assert RAM(26269) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26269))))  severity failure;
	assert RAM(26270) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(26270))))  severity failure;
	assert RAM(26271) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26271))))  severity failure;
	assert RAM(26272) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26272))))  severity failure;
	assert RAM(26273) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(26273))))  severity failure;
	assert RAM(26274) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(26274))))  severity failure;
	assert RAM(26275) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(26275))))  severity failure;
	assert RAM(26276) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(26276))))  severity failure;
	assert RAM(26277) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(26277))))  severity failure;
	assert RAM(26278) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(26278))))  severity failure;
	assert RAM(26279) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(26279))))  severity failure;
	assert RAM(26280) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(26280))))  severity failure;
	assert RAM(26281) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(26281))))  severity failure;
	assert RAM(26282) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(26282))))  severity failure;
	assert RAM(26283) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(26283))))  severity failure;
	assert RAM(26284) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(26284))))  severity failure;
	assert RAM(26285) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(26285))))  severity failure;
	assert RAM(26286) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(26286))))  severity failure;
	assert RAM(26287) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(26287))))  severity failure;
	assert RAM(26288) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26288))))  severity failure;
	assert RAM(26289) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(26289))))  severity failure;
	assert RAM(26290) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(26290))))  severity failure;
	assert RAM(26291) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(26291))))  severity failure;
	assert RAM(26292) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26292))))  severity failure;
	assert RAM(26293) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(26293))))  severity failure;
	assert RAM(26294) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(26294))))  severity failure;
	assert RAM(26295) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26295))))  severity failure;
	assert RAM(26296) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(26296))))  severity failure;
	assert RAM(26297) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(26297))))  severity failure;
	assert RAM(26298) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(26298))))  severity failure;
	assert RAM(26299) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(26299))))  severity failure;
	assert RAM(26300) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26300))))  severity failure;
	assert RAM(26301) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26301))))  severity failure;
	assert RAM(26302) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26302))))  severity failure;
	assert RAM(26303) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(26303))))  severity failure;
	assert RAM(26304) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(26304))))  severity failure;
	assert RAM(26305) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26305))))  severity failure;
	assert RAM(26306) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26306))))  severity failure;
	assert RAM(26307) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26307))))  severity failure;
	assert RAM(26308) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(26308))))  severity failure;
	assert RAM(26309) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(26309))))  severity failure;
	assert RAM(26310) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26310))))  severity failure;
	assert RAM(26311) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(26311))))  severity failure;
	assert RAM(26312) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(26312))))  severity failure;
	assert RAM(26313) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(26313))))  severity failure;
	assert RAM(26314) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(26314))))  severity failure;
	assert RAM(26315) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(26315))))  severity failure;
	assert RAM(26316) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26316))))  severity failure;
	assert RAM(26317) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(26317))))  severity failure;
	assert RAM(26318) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26318))))  severity failure;
	assert RAM(26319) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(26319))))  severity failure;
	assert RAM(26320) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26320))))  severity failure;
	assert RAM(26321) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26321))))  severity failure;
	assert RAM(26322) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(26322))))  severity failure;
	assert RAM(26323) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(26323))))  severity failure;
	assert RAM(26324) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26324))))  severity failure;
	assert RAM(26325) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26325))))  severity failure;
	assert RAM(26326) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(26326))))  severity failure;
	assert RAM(26327) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(26327))))  severity failure;
	assert RAM(26328) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(26328))))  severity failure;
	assert RAM(26329) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(26329))))  severity failure;
	assert RAM(26330) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(26330))))  severity failure;
	assert RAM(26331) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(26331))))  severity failure;
	assert RAM(26332) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(26332))))  severity failure;
	assert RAM(26333) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(26333))))  severity failure;
	assert RAM(26334) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(26334))))  severity failure;
	assert RAM(26335) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26335))))  severity failure;
	assert RAM(26336) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26336))))  severity failure;
	assert RAM(26337) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(26337))))  severity failure;
	assert RAM(26338) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26338))))  severity failure;
	assert RAM(26339) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(26339))))  severity failure;
	assert RAM(26340) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(26340))))  severity failure;
	assert RAM(26341) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26341))))  severity failure;
	assert RAM(26342) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(26342))))  severity failure;
	assert RAM(26343) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26343))))  severity failure;
	assert RAM(26344) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(26344))))  severity failure;
	assert RAM(26345) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(26345))))  severity failure;
	assert RAM(26346) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26346))))  severity failure;
	assert RAM(26347) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(26347))))  severity failure;
	assert RAM(26348) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(26348))))  severity failure;
	assert RAM(26349) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26349))))  severity failure;
	assert RAM(26350) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(26350))))  severity failure;
	assert RAM(26351) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(26351))))  severity failure;
	assert RAM(26352) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(26352))))  severity failure;
	assert RAM(26353) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26353))))  severity failure;
	assert RAM(26354) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26354))))  severity failure;
	assert RAM(26355) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(26355))))  severity failure;
	assert RAM(26356) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26356))))  severity failure;
	assert RAM(26357) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26357))))  severity failure;
	assert RAM(26358) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(26358))))  severity failure;
	assert RAM(26359) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26359))))  severity failure;
	assert RAM(26360) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26360))))  severity failure;
	assert RAM(26361) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26361))))  severity failure;
	assert RAM(26362) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(26362))))  severity failure;
	assert RAM(26363) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(26363))))  severity failure;
	assert RAM(26364) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26364))))  severity failure;
	assert RAM(26365) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(26365))))  severity failure;
	assert RAM(26366) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(26366))))  severity failure;
	assert RAM(26367) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(26367))))  severity failure;
	assert RAM(26368) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(26368))))  severity failure;
	assert RAM(26369) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26369))))  severity failure;
	assert RAM(26370) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(26370))))  severity failure;
	assert RAM(26371) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(26371))))  severity failure;
	assert RAM(26372) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(26372))))  severity failure;
	assert RAM(26373) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26373))))  severity failure;
	assert RAM(26374) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26374))))  severity failure;
	assert RAM(26375) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(26375))))  severity failure;
	assert RAM(26376) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(26376))))  severity failure;
	assert RAM(26377) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(26377))))  severity failure;
	assert RAM(26378) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(26378))))  severity failure;
	assert RAM(26379) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26379))))  severity failure;
	assert RAM(26380) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26380))))  severity failure;
	assert RAM(26381) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(26381))))  severity failure;
	assert RAM(26382) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(26382))))  severity failure;
	assert RAM(26383) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(26383))))  severity failure;
	assert RAM(26384) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26384))))  severity failure;
	assert RAM(26385) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(26385))))  severity failure;
	assert RAM(26386) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(26386))))  severity failure;
	assert RAM(26387) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(26387))))  severity failure;
	assert RAM(26388) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(26388))))  severity failure;
	assert RAM(26389) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(26389))))  severity failure;
	assert RAM(26390) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(26390))))  severity failure;
	assert RAM(26391) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(26391))))  severity failure;
	assert RAM(26392) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(26392))))  severity failure;
	assert RAM(26393) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26393))))  severity failure;
	assert RAM(26394) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(26394))))  severity failure;
	assert RAM(26395) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26395))))  severity failure;
	assert RAM(26396) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(26396))))  severity failure;
	assert RAM(26397) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(26397))))  severity failure;
	assert RAM(26398) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(26398))))  severity failure;
	assert RAM(26399) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(26399))))  severity failure;
	assert RAM(26400) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(26400))))  severity failure;
	assert RAM(26401) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(26401))))  severity failure;
	assert RAM(26402) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(26402))))  severity failure;
	assert RAM(26403) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(26403))))  severity failure;
	assert RAM(26404) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(26404))))  severity failure;
	assert RAM(26405) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(26405))))  severity failure;
	assert RAM(26406) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(26406))))  severity failure;
	assert RAM(26407) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26407))))  severity failure;
	assert RAM(26408) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26408))))  severity failure;
	assert RAM(26409) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(26409))))  severity failure;
	assert RAM(26410) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26410))))  severity failure;
	assert RAM(26411) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(26411))))  severity failure;
	assert RAM(26412) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(26412))))  severity failure;
	assert RAM(26413) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(26413))))  severity failure;
	assert RAM(26414) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(26414))))  severity failure;
	assert RAM(26415) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(26415))))  severity failure;
	assert RAM(26416) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26416))))  severity failure;
	assert RAM(26417) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(26417))))  severity failure;
	assert RAM(26418) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(26418))))  severity failure;
	assert RAM(26419) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26419))))  severity failure;
	assert RAM(26420) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(26420))))  severity failure;
	assert RAM(26421) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(26421))))  severity failure;
	assert RAM(26422) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26422))))  severity failure;
	assert RAM(26423) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26423))))  severity failure;
	assert RAM(26424) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(26424))))  severity failure;
	assert RAM(26425) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26425))))  severity failure;
	assert RAM(26426) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(26426))))  severity failure;
	assert RAM(26427) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(26427))))  severity failure;
	assert RAM(26428) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(26428))))  severity failure;
	assert RAM(26429) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26429))))  severity failure;
	assert RAM(26430) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(26430))))  severity failure;
	assert RAM(26431) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26431))))  severity failure;
	assert RAM(26432) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26432))))  severity failure;
	assert RAM(26433) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(26433))))  severity failure;
	assert RAM(26434) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(26434))))  severity failure;
	assert RAM(26435) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(26435))))  severity failure;
	assert RAM(26436) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26436))))  severity failure;
	assert RAM(26437) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26437))))  severity failure;
	assert RAM(26438) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(26438))))  severity failure;
	assert RAM(26439) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(26439))))  severity failure;
	assert RAM(26440) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(26440))))  severity failure;
	assert RAM(26441) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(26441))))  severity failure;
	assert RAM(26442) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26442))))  severity failure;
	assert RAM(26443) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(26443))))  severity failure;
	assert RAM(26444) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26444))))  severity failure;
	assert RAM(26445) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(26445))))  severity failure;
	assert RAM(26446) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(26446))))  severity failure;
	assert RAM(26447) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(26447))))  severity failure;
	assert RAM(26448) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26448))))  severity failure;
	assert RAM(26449) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26449))))  severity failure;
	assert RAM(26450) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26450))))  severity failure;
	assert RAM(26451) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(26451))))  severity failure;
	assert RAM(26452) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26452))))  severity failure;
	assert RAM(26453) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(26453))))  severity failure;
	assert RAM(26454) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(26454))))  severity failure;
	assert RAM(26455) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26455))))  severity failure;
	assert RAM(26456) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(26456))))  severity failure;
	assert RAM(26457) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(26457))))  severity failure;
	assert RAM(26458) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26458))))  severity failure;
	assert RAM(26459) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(26459))))  severity failure;
	assert RAM(26460) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26460))))  severity failure;
	assert RAM(26461) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(26461))))  severity failure;
	assert RAM(26462) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26462))))  severity failure;
	assert RAM(26463) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(26463))))  severity failure;
	assert RAM(26464) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(26464))))  severity failure;
	assert RAM(26465) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26465))))  severity failure;
	assert RAM(26466) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26466))))  severity failure;
	assert RAM(26467) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26467))))  severity failure;
	assert RAM(26468) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26468))))  severity failure;
	assert RAM(26469) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(26469))))  severity failure;
	assert RAM(26470) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(26470))))  severity failure;
	assert RAM(26471) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(26471))))  severity failure;
	assert RAM(26472) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(26472))))  severity failure;
	assert RAM(26473) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(26473))))  severity failure;
	assert RAM(26474) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(26474))))  severity failure;
	assert RAM(26475) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(26475))))  severity failure;
	assert RAM(26476) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(26476))))  severity failure;
	assert RAM(26477) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26477))))  severity failure;
	assert RAM(26478) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(26478))))  severity failure;
	assert RAM(26479) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26479))))  severity failure;
	assert RAM(26480) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(26480))))  severity failure;
	assert RAM(26481) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(26481))))  severity failure;
	assert RAM(26482) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(26482))))  severity failure;
	assert RAM(26483) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(26483))))  severity failure;
	assert RAM(26484) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26484))))  severity failure;
	assert RAM(26485) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(26485))))  severity failure;
	assert RAM(26486) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26486))))  severity failure;
	assert RAM(26487) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(26487))))  severity failure;
	assert RAM(26488) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(26488))))  severity failure;
	assert RAM(26489) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(26489))))  severity failure;
	assert RAM(26490) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(26490))))  severity failure;
	assert RAM(26491) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(26491))))  severity failure;
	assert RAM(26492) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26492))))  severity failure;
	assert RAM(26493) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(26493))))  severity failure;
	assert RAM(26494) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(26494))))  severity failure;
	assert RAM(26495) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(26495))))  severity failure;
	assert RAM(26496) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(26496))))  severity failure;
	assert RAM(26497) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26497))))  severity failure;
	assert RAM(26498) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(26498))))  severity failure;
	assert RAM(26499) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26499))))  severity failure;
	assert RAM(26500) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(26500))))  severity failure;
	assert RAM(26501) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(26501))))  severity failure;
	assert RAM(26502) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26502))))  severity failure;
	assert RAM(26503) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(26503))))  severity failure;
	assert RAM(26504) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(26504))))  severity failure;
	assert RAM(26505) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(26505))))  severity failure;
	assert RAM(26506) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(26506))))  severity failure;
	assert RAM(26507) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26507))))  severity failure;
	assert RAM(26508) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(26508))))  severity failure;
	assert RAM(26509) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(26509))))  severity failure;
	assert RAM(26510) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26510))))  severity failure;
	assert RAM(26511) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26511))))  severity failure;
	assert RAM(26512) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(26512))))  severity failure;
	assert RAM(26513) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(26513))))  severity failure;
	assert RAM(26514) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(26514))))  severity failure;
	assert RAM(26515) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(26515))))  severity failure;
	assert RAM(26516) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26516))))  severity failure;
	assert RAM(26517) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26517))))  severity failure;
	assert RAM(26518) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26518))))  severity failure;
	assert RAM(26519) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(26519))))  severity failure;
	assert RAM(26520) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26520))))  severity failure;
	assert RAM(26521) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26521))))  severity failure;
	assert RAM(26522) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(26522))))  severity failure;
	assert RAM(26523) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(26523))))  severity failure;
	assert RAM(26524) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26524))))  severity failure;
	assert RAM(26525) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26525))))  severity failure;
	assert RAM(26526) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26526))))  severity failure;
	assert RAM(26527) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26527))))  severity failure;
	assert RAM(26528) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(26528))))  severity failure;
	assert RAM(26529) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(26529))))  severity failure;
	assert RAM(26530) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26530))))  severity failure;
	assert RAM(26531) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(26531))))  severity failure;
	assert RAM(26532) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(26532))))  severity failure;
	assert RAM(26533) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(26533))))  severity failure;
	assert RAM(26534) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(26534))))  severity failure;
	assert RAM(26535) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(26535))))  severity failure;
	assert RAM(26536) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(26536))))  severity failure;
	assert RAM(26537) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(26537))))  severity failure;
	assert RAM(26538) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(26538))))  severity failure;
	assert RAM(26539) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(26539))))  severity failure;
	assert RAM(26540) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(26540))))  severity failure;
	assert RAM(26541) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(26541))))  severity failure;
	assert RAM(26542) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(26542))))  severity failure;
	assert RAM(26543) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(26543))))  severity failure;
	assert RAM(26544) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(26544))))  severity failure;
	assert RAM(26545) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(26545))))  severity failure;
	assert RAM(26546) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26546))))  severity failure;
	assert RAM(26547) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26547))))  severity failure;
	assert RAM(26548) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(26548))))  severity failure;
	assert RAM(26549) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(26549))))  severity failure;
	assert RAM(26550) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(26550))))  severity failure;
	assert RAM(26551) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(26551))))  severity failure;
	assert RAM(26552) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26552))))  severity failure;
	assert RAM(26553) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(26553))))  severity failure;
	assert RAM(26554) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(26554))))  severity failure;
	assert RAM(26555) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(26555))))  severity failure;
	assert RAM(26556) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26556))))  severity failure;
	assert RAM(26557) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(26557))))  severity failure;
	assert RAM(26558) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26558))))  severity failure;
	assert RAM(26559) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(26559))))  severity failure;
	assert RAM(26560) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(26560))))  severity failure;
	assert RAM(26561) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26561))))  severity failure;
	assert RAM(26562) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(26562))))  severity failure;
	assert RAM(26563) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26563))))  severity failure;
	assert RAM(26564) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(26564))))  severity failure;
	assert RAM(26565) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(26565))))  severity failure;
	assert RAM(26566) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(26566))))  severity failure;
	assert RAM(26567) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26567))))  severity failure;
	assert RAM(26568) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26568))))  severity failure;
	assert RAM(26569) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(26569))))  severity failure;
	assert RAM(26570) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(26570))))  severity failure;
	assert RAM(26571) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26571))))  severity failure;
	assert RAM(26572) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(26572))))  severity failure;
	assert RAM(26573) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26573))))  severity failure;
	assert RAM(26574) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(26574))))  severity failure;
	assert RAM(26575) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(26575))))  severity failure;
	assert RAM(26576) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(26576))))  severity failure;
	assert RAM(26577) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(26577))))  severity failure;
	assert RAM(26578) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(26578))))  severity failure;
	assert RAM(26579) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(26579))))  severity failure;
	assert RAM(26580) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26580))))  severity failure;
	assert RAM(26581) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26581))))  severity failure;
	assert RAM(26582) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26582))))  severity failure;
	assert RAM(26583) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(26583))))  severity failure;
	assert RAM(26584) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26584))))  severity failure;
	assert RAM(26585) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(26585))))  severity failure;
	assert RAM(26586) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(26586))))  severity failure;
	assert RAM(26587) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(26587))))  severity failure;
	assert RAM(26588) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26588))))  severity failure;
	assert RAM(26589) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(26589))))  severity failure;
	assert RAM(26590) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26590))))  severity failure;
	assert RAM(26591) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(26591))))  severity failure;
	assert RAM(26592) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(26592))))  severity failure;
	assert RAM(26593) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(26593))))  severity failure;
	assert RAM(26594) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(26594))))  severity failure;
	assert RAM(26595) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26595))))  severity failure;
	assert RAM(26596) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26596))))  severity failure;
	assert RAM(26597) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(26597))))  severity failure;
	assert RAM(26598) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(26598))))  severity failure;
	assert RAM(26599) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(26599))))  severity failure;
	assert RAM(26600) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26600))))  severity failure;
	assert RAM(26601) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(26601))))  severity failure;
	assert RAM(26602) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(26602))))  severity failure;
	assert RAM(26603) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(26603))))  severity failure;
	assert RAM(26604) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(26604))))  severity failure;
	assert RAM(26605) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(26605))))  severity failure;
	assert RAM(26606) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26606))))  severity failure;
	assert RAM(26607) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(26607))))  severity failure;
	assert RAM(26608) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(26608))))  severity failure;
	assert RAM(26609) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26609))))  severity failure;
	assert RAM(26610) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(26610))))  severity failure;
	assert RAM(26611) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(26611))))  severity failure;
	assert RAM(26612) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(26612))))  severity failure;
	assert RAM(26613) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(26613))))  severity failure;
	assert RAM(26614) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(26614))))  severity failure;
	assert RAM(26615) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26615))))  severity failure;
	assert RAM(26616) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(26616))))  severity failure;
	assert RAM(26617) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(26617))))  severity failure;
	assert RAM(26618) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26618))))  severity failure;
	assert RAM(26619) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(26619))))  severity failure;
	assert RAM(26620) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26620))))  severity failure;
	assert RAM(26621) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26621))))  severity failure;
	assert RAM(26622) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(26622))))  severity failure;
	assert RAM(26623) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26623))))  severity failure;
	assert RAM(26624) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(26624))))  severity failure;
	assert RAM(26625) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(26625))))  severity failure;
	assert RAM(26626) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26626))))  severity failure;
	assert RAM(26627) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(26627))))  severity failure;
	assert RAM(26628) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(26628))))  severity failure;
	assert RAM(26629) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26629))))  severity failure;
	assert RAM(26630) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(26630))))  severity failure;
	assert RAM(26631) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(26631))))  severity failure;
	assert RAM(26632) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(26632))))  severity failure;
	assert RAM(26633) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(26633))))  severity failure;
	assert RAM(26634) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(26634))))  severity failure;
	assert RAM(26635) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(26635))))  severity failure;
	assert RAM(26636) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(26636))))  severity failure;
	assert RAM(26637) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(26637))))  severity failure;
	assert RAM(26638) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(26638))))  severity failure;
	assert RAM(26639) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26639))))  severity failure;
	assert RAM(26640) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26640))))  severity failure;
	assert RAM(26641) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(26641))))  severity failure;
	assert RAM(26642) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(26642))))  severity failure;
	assert RAM(26643) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(26643))))  severity failure;
	assert RAM(26644) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26644))))  severity failure;
	assert RAM(26645) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(26645))))  severity failure;
	assert RAM(26646) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26646))))  severity failure;
	assert RAM(26647) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(26647))))  severity failure;
	assert RAM(26648) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(26648))))  severity failure;
	assert RAM(26649) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26649))))  severity failure;
	assert RAM(26650) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(26650))))  severity failure;
	assert RAM(26651) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(26651))))  severity failure;
	assert RAM(26652) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(26652))))  severity failure;
	assert RAM(26653) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(26653))))  severity failure;
	assert RAM(26654) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(26654))))  severity failure;
	assert RAM(26655) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(26655))))  severity failure;
	assert RAM(26656) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(26656))))  severity failure;
	assert RAM(26657) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26657))))  severity failure;
	assert RAM(26658) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26658))))  severity failure;
	assert RAM(26659) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(26659))))  severity failure;
	assert RAM(26660) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(26660))))  severity failure;
	assert RAM(26661) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(26661))))  severity failure;
	assert RAM(26662) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(26662))))  severity failure;
	assert RAM(26663) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(26663))))  severity failure;
	assert RAM(26664) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(26664))))  severity failure;
	assert RAM(26665) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(26665))))  severity failure;
	assert RAM(26666) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(26666))))  severity failure;
	assert RAM(26667) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(26667))))  severity failure;
	assert RAM(26668) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(26668))))  severity failure;
	assert RAM(26669) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(26669))))  severity failure;
	assert RAM(26670) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(26670))))  severity failure;
	assert RAM(26671) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(26671))))  severity failure;
	assert RAM(26672) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26672))))  severity failure;
	assert RAM(26673) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(26673))))  severity failure;
	assert RAM(26674) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(26674))))  severity failure;
	assert RAM(26675) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(26675))))  severity failure;
	assert RAM(26676) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26676))))  severity failure;
	assert RAM(26677) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(26677))))  severity failure;
	assert RAM(26678) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(26678))))  severity failure;
	assert RAM(26679) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26679))))  severity failure;
	assert RAM(26680) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26680))))  severity failure;
	assert RAM(26681) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(26681))))  severity failure;
	assert RAM(26682) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(26682))))  severity failure;
	assert RAM(26683) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(26683))))  severity failure;
	assert RAM(26684) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(26684))))  severity failure;
	assert RAM(26685) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26685))))  severity failure;
	assert RAM(26686) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26686))))  severity failure;
	assert RAM(26687) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(26687))))  severity failure;
	assert RAM(26688) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(26688))))  severity failure;
	assert RAM(26689) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(26689))))  severity failure;
	assert RAM(26690) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26690))))  severity failure;
	assert RAM(26691) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(26691))))  severity failure;
	assert RAM(26692) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(26692))))  severity failure;
	assert RAM(26693) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26693))))  severity failure;
	assert RAM(26694) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26694))))  severity failure;
	assert RAM(26695) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(26695))))  severity failure;
	assert RAM(26696) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26696))))  severity failure;
	assert RAM(26697) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(26697))))  severity failure;
	assert RAM(26698) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(26698))))  severity failure;
	assert RAM(26699) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(26699))))  severity failure;
	assert RAM(26700) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(26700))))  severity failure;
	assert RAM(26701) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(26701))))  severity failure;
	assert RAM(26702) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(26702))))  severity failure;
	assert RAM(26703) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(26703))))  severity failure;
	assert RAM(26704) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(26704))))  severity failure;
	assert RAM(26705) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(26705))))  severity failure;
	assert RAM(26706) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26706))))  severity failure;
	assert RAM(26707) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(26707))))  severity failure;
	assert RAM(26708) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(26708))))  severity failure;
	assert RAM(26709) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26709))))  severity failure;
	assert RAM(26710) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26710))))  severity failure;
	assert RAM(26711) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(26711))))  severity failure;
	assert RAM(26712) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(26712))))  severity failure;
	assert RAM(26713) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(26713))))  severity failure;
	assert RAM(26714) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26714))))  severity failure;
	assert RAM(26715) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(26715))))  severity failure;
	assert RAM(26716) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26716))))  severity failure;
	assert RAM(26717) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26717))))  severity failure;
	assert RAM(26718) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26718))))  severity failure;
	assert RAM(26719) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(26719))))  severity failure;
	assert RAM(26720) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(26720))))  severity failure;
	assert RAM(26721) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26721))))  severity failure;
	assert RAM(26722) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(26722))))  severity failure;
	assert RAM(26723) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26723))))  severity failure;
	assert RAM(26724) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(26724))))  severity failure;
	assert RAM(26725) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26725))))  severity failure;
	assert RAM(26726) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26726))))  severity failure;
	assert RAM(26727) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(26727))))  severity failure;
	assert RAM(26728) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26728))))  severity failure;
	assert RAM(26729) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(26729))))  severity failure;
	assert RAM(26730) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(26730))))  severity failure;
	assert RAM(26731) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(26731))))  severity failure;
	assert RAM(26732) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(26732))))  severity failure;
	assert RAM(26733) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26733))))  severity failure;
	assert RAM(26734) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26734))))  severity failure;
	assert RAM(26735) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26735))))  severity failure;
	assert RAM(26736) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(26736))))  severity failure;
	assert RAM(26737) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(26737))))  severity failure;
	assert RAM(26738) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(26738))))  severity failure;
	assert RAM(26739) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(26739))))  severity failure;
	assert RAM(26740) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(26740))))  severity failure;
	assert RAM(26741) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(26741))))  severity failure;
	assert RAM(26742) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(26742))))  severity failure;
	assert RAM(26743) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(26743))))  severity failure;
	assert RAM(26744) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26744))))  severity failure;
	assert RAM(26745) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(26745))))  severity failure;
	assert RAM(26746) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(26746))))  severity failure;
	assert RAM(26747) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(26747))))  severity failure;
	assert RAM(26748) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(26748))))  severity failure;
	assert RAM(26749) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(26749))))  severity failure;
	assert RAM(26750) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(26750))))  severity failure;
	assert RAM(26751) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(26751))))  severity failure;
	assert RAM(26752) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(26752))))  severity failure;
	assert RAM(26753) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26753))))  severity failure;
	assert RAM(26754) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(26754))))  severity failure;
	assert RAM(26755) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(26755))))  severity failure;
	assert RAM(26756) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26756))))  severity failure;
	assert RAM(26757) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(26757))))  severity failure;
	assert RAM(26758) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(26758))))  severity failure;
	assert RAM(26759) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(26759))))  severity failure;
	assert RAM(26760) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(26760))))  severity failure;
	assert RAM(26761) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(26761))))  severity failure;
	assert RAM(26762) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(26762))))  severity failure;
	assert RAM(26763) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26763))))  severity failure;
	assert RAM(26764) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(26764))))  severity failure;
	assert RAM(26765) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26765))))  severity failure;
	assert RAM(26766) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26766))))  severity failure;
	assert RAM(26767) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(26767))))  severity failure;
	assert RAM(26768) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(26768))))  severity failure;
	assert RAM(26769) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(26769))))  severity failure;
	assert RAM(26770) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26770))))  severity failure;
	assert RAM(26771) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26771))))  severity failure;
	assert RAM(26772) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(26772))))  severity failure;
	assert RAM(26773) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(26773))))  severity failure;
	assert RAM(26774) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26774))))  severity failure;
	assert RAM(26775) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26775))))  severity failure;
	assert RAM(26776) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(26776))))  severity failure;
	assert RAM(26777) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(26777))))  severity failure;
	assert RAM(26778) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(26778))))  severity failure;
	assert RAM(26779) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(26779))))  severity failure;
	assert RAM(26780) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(26780))))  severity failure;
	assert RAM(26781) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26781))))  severity failure;
	assert RAM(26782) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(26782))))  severity failure;
	assert RAM(26783) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(26783))))  severity failure;
	assert RAM(26784) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26784))))  severity failure;
	assert RAM(26785) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(26785))))  severity failure;
	assert RAM(26786) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(26786))))  severity failure;
	assert RAM(26787) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26787))))  severity failure;
	assert RAM(26788) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26788))))  severity failure;
	assert RAM(26789) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(26789))))  severity failure;
	assert RAM(26790) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(26790))))  severity failure;
	assert RAM(26791) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(26791))))  severity failure;
	assert RAM(26792) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(26792))))  severity failure;
	assert RAM(26793) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(26793))))  severity failure;
	assert RAM(26794) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(26794))))  severity failure;
	assert RAM(26795) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(26795))))  severity failure;
	assert RAM(26796) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(26796))))  severity failure;
	assert RAM(26797) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(26797))))  severity failure;
	assert RAM(26798) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(26798))))  severity failure;
	assert RAM(26799) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26799))))  severity failure;
	assert RAM(26800) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(26800))))  severity failure;
	assert RAM(26801) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(26801))))  severity failure;
	assert RAM(26802) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26802))))  severity failure;
	assert RAM(26803) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(26803))))  severity failure;
	assert RAM(26804) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26804))))  severity failure;
	assert RAM(26805) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(26805))))  severity failure;
	assert RAM(26806) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(26806))))  severity failure;
	assert RAM(26807) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(26807))))  severity failure;
	assert RAM(26808) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(26808))))  severity failure;
	assert RAM(26809) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26809))))  severity failure;
	assert RAM(26810) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(26810))))  severity failure;
	assert RAM(26811) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(26811))))  severity failure;
	assert RAM(26812) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(26812))))  severity failure;
	assert RAM(26813) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26813))))  severity failure;
	assert RAM(26814) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(26814))))  severity failure;
	assert RAM(26815) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26815))))  severity failure;
	assert RAM(26816) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(26816))))  severity failure;
	assert RAM(26817) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(26817))))  severity failure;
	assert RAM(26818) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(26818))))  severity failure;
	assert RAM(26819) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26819))))  severity failure;
	assert RAM(26820) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(26820))))  severity failure;
	assert RAM(26821) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(26821))))  severity failure;
	assert RAM(26822) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(26822))))  severity failure;
	assert RAM(26823) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(26823))))  severity failure;
	assert RAM(26824) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26824))))  severity failure;
	assert RAM(26825) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(26825))))  severity failure;
	assert RAM(26826) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(26826))))  severity failure;
	assert RAM(26827) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(26827))))  severity failure;
	assert RAM(26828) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(26828))))  severity failure;
	assert RAM(26829) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26829))))  severity failure;
	assert RAM(26830) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(26830))))  severity failure;
	assert RAM(26831) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(26831))))  severity failure;
	assert RAM(26832) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26832))))  severity failure;
	assert RAM(26833) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(26833))))  severity failure;
	assert RAM(26834) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(26834))))  severity failure;
	assert RAM(26835) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(26835))))  severity failure;
	assert RAM(26836) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26836))))  severity failure;
	assert RAM(26837) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(26837))))  severity failure;
	assert RAM(26838) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(26838))))  severity failure;
	assert RAM(26839) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(26839))))  severity failure;
	assert RAM(26840) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26840))))  severity failure;
	assert RAM(26841) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(26841))))  severity failure;
	assert RAM(26842) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26842))))  severity failure;
	assert RAM(26843) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(26843))))  severity failure;
	assert RAM(26844) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(26844))))  severity failure;
	assert RAM(26845) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(26845))))  severity failure;
	assert RAM(26846) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(26846))))  severity failure;
	assert RAM(26847) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(26847))))  severity failure;
	assert RAM(26848) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(26848))))  severity failure;
	assert RAM(26849) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(26849))))  severity failure;
	assert RAM(26850) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(26850))))  severity failure;
	assert RAM(26851) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(26851))))  severity failure;
	assert RAM(26852) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(26852))))  severity failure;
	assert RAM(26853) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(26853))))  severity failure;
	assert RAM(26854) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(26854))))  severity failure;
	assert RAM(26855) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(26855))))  severity failure;
	assert RAM(26856) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26856))))  severity failure;
	assert RAM(26857) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(26857))))  severity failure;
	assert RAM(26858) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(26858))))  severity failure;
	assert RAM(26859) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(26859))))  severity failure;
	assert RAM(26860) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(26860))))  severity failure;
	assert RAM(26861) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26861))))  severity failure;
	assert RAM(26862) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(26862))))  severity failure;
	assert RAM(26863) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(26863))))  severity failure;
	assert RAM(26864) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(26864))))  severity failure;
	assert RAM(26865) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(26865))))  severity failure;
	assert RAM(26866) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(26866))))  severity failure;
	assert RAM(26867) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(26867))))  severity failure;
	assert RAM(26868) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(26868))))  severity failure;
	assert RAM(26869) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(26869))))  severity failure;
	assert RAM(26870) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(26870))))  severity failure;
	assert RAM(26871) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(26871))))  severity failure;
	assert RAM(26872) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(26872))))  severity failure;
	assert RAM(26873) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(26873))))  severity failure;
	assert RAM(26874) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(26874))))  severity failure;
	assert RAM(26875) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26875))))  severity failure;
	assert RAM(26876) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(26876))))  severity failure;
	assert RAM(26877) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(26877))))  severity failure;
	assert RAM(26878) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(26878))))  severity failure;
	assert RAM(26879) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(26879))))  severity failure;
	assert RAM(26880) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(26880))))  severity failure;
	assert RAM(26881) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(26881))))  severity failure;
	assert RAM(26882) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(26882))))  severity failure;
	assert RAM(26883) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(26883))))  severity failure;
	assert RAM(26884) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(26884))))  severity failure;
	assert RAM(26885) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(26885))))  severity failure;
	assert RAM(26886) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(26886))))  severity failure;
	assert RAM(26887) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(26887))))  severity failure;
	assert RAM(26888) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(26888))))  severity failure;
	assert RAM(26889) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(26889))))  severity failure;
	assert RAM(26890) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26890))))  severity failure;
	assert RAM(26891) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(26891))))  severity failure;
	assert RAM(26892) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(26892))))  severity failure;
	assert RAM(26893) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(26893))))  severity failure;
	assert RAM(26894) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(26894))))  severity failure;
	assert RAM(26895) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(26895))))  severity failure;
	assert RAM(26896) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26896))))  severity failure;
	assert RAM(26897) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(26897))))  severity failure;
	assert RAM(26898) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(26898))))  severity failure;
	assert RAM(26899) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(26899))))  severity failure;
	assert RAM(26900) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(26900))))  severity failure;
	assert RAM(26901) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(26901))))  severity failure;
	assert RAM(26902) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26902))))  severity failure;
	assert RAM(26903) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26903))))  severity failure;
	assert RAM(26904) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(26904))))  severity failure;
	assert RAM(26905) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(26905))))  severity failure;
	assert RAM(26906) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(26906))))  severity failure;
	assert RAM(26907) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26907))))  severity failure;
	assert RAM(26908) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(26908))))  severity failure;
	assert RAM(26909) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(26909))))  severity failure;
	assert RAM(26910) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(26910))))  severity failure;
	assert RAM(26911) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(26911))))  severity failure;
	assert RAM(26912) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(26912))))  severity failure;
	assert RAM(26913) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(26913))))  severity failure;
	assert RAM(26914) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(26914))))  severity failure;
	assert RAM(26915) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(26915))))  severity failure;
	assert RAM(26916) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(26916))))  severity failure;
	assert RAM(26917) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(26917))))  severity failure;
	assert RAM(26918) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(26918))))  severity failure;
	assert RAM(26919) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26919))))  severity failure;
	assert RAM(26920) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(26920))))  severity failure;
	assert RAM(26921) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(26921))))  severity failure;
	assert RAM(26922) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(26922))))  severity failure;
	assert RAM(26923) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(26923))))  severity failure;
	assert RAM(26924) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(26924))))  severity failure;
	assert RAM(26925) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26925))))  severity failure;
	assert RAM(26926) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(26926))))  severity failure;
	assert RAM(26927) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(26927))))  severity failure;
	assert RAM(26928) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26928))))  severity failure;
	assert RAM(26929) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(26929))))  severity failure;
	assert RAM(26930) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(26930))))  severity failure;
	assert RAM(26931) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(26931))))  severity failure;
	assert RAM(26932) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(26932))))  severity failure;
	assert RAM(26933) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(26933))))  severity failure;
	assert RAM(26934) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(26934))))  severity failure;
	assert RAM(26935) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(26935))))  severity failure;
	assert RAM(26936) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26936))))  severity failure;
	assert RAM(26937) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(26937))))  severity failure;
	assert RAM(26938) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(26938))))  severity failure;
	assert RAM(26939) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(26939))))  severity failure;
	assert RAM(26940) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(26940))))  severity failure;
	assert RAM(26941) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(26941))))  severity failure;
	assert RAM(26942) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(26942))))  severity failure;
	assert RAM(26943) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(26943))))  severity failure;
	assert RAM(26944) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26944))))  severity failure;
	assert RAM(26945) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(26945))))  severity failure;
	assert RAM(26946) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(26946))))  severity failure;
	assert RAM(26947) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(26947))))  severity failure;
	assert RAM(26948) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(26948))))  severity failure;
	assert RAM(26949) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(26949))))  severity failure;
	assert RAM(26950) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(26950))))  severity failure;
	assert RAM(26951) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(26951))))  severity failure;
	assert RAM(26952) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(26952))))  severity failure;
	assert RAM(26953) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26953))))  severity failure;
	assert RAM(26954) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(26954))))  severity failure;
	assert RAM(26955) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(26955))))  severity failure;
	assert RAM(26956) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26956))))  severity failure;
	assert RAM(26957) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(26957))))  severity failure;
	assert RAM(26958) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(26958))))  severity failure;
	assert RAM(26959) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(26959))))  severity failure;
	assert RAM(26960) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(26960))))  severity failure;
	assert RAM(26961) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(26961))))  severity failure;
	assert RAM(26962) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(26962))))  severity failure;
	assert RAM(26963) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(26963))))  severity failure;
	assert RAM(26964) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(26964))))  severity failure;
	assert RAM(26965) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(26965))))  severity failure;
	assert RAM(26966) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(26966))))  severity failure;
	assert RAM(26967) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(26967))))  severity failure;
	assert RAM(26968) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(26968))))  severity failure;
	assert RAM(26969) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(26969))))  severity failure;
	assert RAM(26970) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(26970))))  severity failure;
	assert RAM(26971) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(26971))))  severity failure;
	assert RAM(26972) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(26972))))  severity failure;
	assert RAM(26973) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(26973))))  severity failure;
	assert RAM(26974) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(26974))))  severity failure;
	assert RAM(26975) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(26975))))  severity failure;
	assert RAM(26976) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(26976))))  severity failure;
	assert RAM(26977) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(26977))))  severity failure;
	assert RAM(26978) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(26978))))  severity failure;
	assert RAM(26979) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(26979))))  severity failure;
	assert RAM(26980) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26980))))  severity failure;
	assert RAM(26981) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(26981))))  severity failure;
	assert RAM(26982) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(26982))))  severity failure;
	assert RAM(26983) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(26983))))  severity failure;
	assert RAM(26984) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(26984))))  severity failure;
	assert RAM(26985) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(26985))))  severity failure;
	assert RAM(26986) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(26986))))  severity failure;
	assert RAM(26987) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(26987))))  severity failure;
	assert RAM(26988) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(26988))))  severity failure;
	assert RAM(26989) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(26989))))  severity failure;
	assert RAM(26990) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(26990))))  severity failure;
	assert RAM(26991) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(26991))))  severity failure;
	assert RAM(26992) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(26992))))  severity failure;
	assert RAM(26993) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(26993))))  severity failure;
	assert RAM(26994) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(26994))))  severity failure;
	assert RAM(26995) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(26995))))  severity failure;
	assert RAM(26996) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(26996))))  severity failure;
	assert RAM(26997) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(26997))))  severity failure;
	assert RAM(26998) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(26998))))  severity failure;
	assert RAM(26999) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(26999))))  severity failure;
	assert RAM(27000) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(27000))))  severity failure;
	assert RAM(27001) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(27001))))  severity failure;
	assert RAM(27002) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27002))))  severity failure;
	assert RAM(27003) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(27003))))  severity failure;
	assert RAM(27004) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27004))))  severity failure;
	assert RAM(27005) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(27005))))  severity failure;
	assert RAM(27006) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27006))))  severity failure;
	assert RAM(27007) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27007))))  severity failure;
	assert RAM(27008) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(27008))))  severity failure;
	assert RAM(27009) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(27009))))  severity failure;
	assert RAM(27010) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(27010))))  severity failure;
	assert RAM(27011) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(27011))))  severity failure;
	assert RAM(27012) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27012))))  severity failure;
	assert RAM(27013) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27013))))  severity failure;
	assert RAM(27014) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27014))))  severity failure;
	assert RAM(27015) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(27015))))  severity failure;
	assert RAM(27016) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27016))))  severity failure;
	assert RAM(27017) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(27017))))  severity failure;
	assert RAM(27018) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27018))))  severity failure;
	assert RAM(27019) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27019))))  severity failure;
	assert RAM(27020) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(27020))))  severity failure;
	assert RAM(27021) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(27021))))  severity failure;
	assert RAM(27022) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27022))))  severity failure;
	assert RAM(27023) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(27023))))  severity failure;
	assert RAM(27024) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(27024))))  severity failure;
	assert RAM(27025) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(27025))))  severity failure;
	assert RAM(27026) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(27026))))  severity failure;
	assert RAM(27027) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(27027))))  severity failure;
	assert RAM(27028) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27028))))  severity failure;
	assert RAM(27029) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(27029))))  severity failure;
	assert RAM(27030) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27030))))  severity failure;
	assert RAM(27031) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(27031))))  severity failure;
	assert RAM(27032) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(27032))))  severity failure;
	assert RAM(27033) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27033))))  severity failure;
	assert RAM(27034) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(27034))))  severity failure;
	assert RAM(27035) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(27035))))  severity failure;
	assert RAM(27036) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27036))))  severity failure;
	assert RAM(27037) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(27037))))  severity failure;
	assert RAM(27038) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27038))))  severity failure;
	assert RAM(27039) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(27039))))  severity failure;
	assert RAM(27040) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(27040))))  severity failure;
	assert RAM(27041) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(27041))))  severity failure;
	assert RAM(27042) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(27042))))  severity failure;
	assert RAM(27043) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(27043))))  severity failure;
	assert RAM(27044) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(27044))))  severity failure;
	assert RAM(27045) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(27045))))  severity failure;
	assert RAM(27046) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27046))))  severity failure;
	assert RAM(27047) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27047))))  severity failure;
	assert RAM(27048) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27048))))  severity failure;
	assert RAM(27049) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(27049))))  severity failure;
	assert RAM(27050) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(27050))))  severity failure;
	assert RAM(27051) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(27051))))  severity failure;
	assert RAM(27052) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(27052))))  severity failure;
	assert RAM(27053) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27053))))  severity failure;
	assert RAM(27054) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(27054))))  severity failure;
	assert RAM(27055) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(27055))))  severity failure;
	assert RAM(27056) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27056))))  severity failure;
	assert RAM(27057) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(27057))))  severity failure;
	assert RAM(27058) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27058))))  severity failure;
	assert RAM(27059) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27059))))  severity failure;
	assert RAM(27060) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27060))))  severity failure;
	assert RAM(27061) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27061))))  severity failure;
	assert RAM(27062) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27062))))  severity failure;
	assert RAM(27063) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(27063))))  severity failure;
	assert RAM(27064) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(27064))))  severity failure;
	assert RAM(27065) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(27065))))  severity failure;
	assert RAM(27066) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(27066))))  severity failure;
	assert RAM(27067) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27067))))  severity failure;
	assert RAM(27068) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(27068))))  severity failure;
	assert RAM(27069) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(27069))))  severity failure;
	assert RAM(27070) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27070))))  severity failure;
	assert RAM(27071) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(27071))))  severity failure;
	assert RAM(27072) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(27072))))  severity failure;
	assert RAM(27073) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(27073))))  severity failure;
	assert RAM(27074) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(27074))))  severity failure;
	assert RAM(27075) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(27075))))  severity failure;
	assert RAM(27076) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27076))))  severity failure;
	assert RAM(27077) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(27077))))  severity failure;
	assert RAM(27078) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27078))))  severity failure;
	assert RAM(27079) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(27079))))  severity failure;
	assert RAM(27080) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27080))))  severity failure;
	assert RAM(27081) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(27081))))  severity failure;
	assert RAM(27082) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27082))))  severity failure;
	assert RAM(27083) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(27083))))  severity failure;
	assert RAM(27084) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(27084))))  severity failure;
	assert RAM(27085) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(27085))))  severity failure;
	assert RAM(27086) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(27086))))  severity failure;
	assert RAM(27087) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27087))))  severity failure;
	assert RAM(27088) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(27088))))  severity failure;
	assert RAM(27089) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27089))))  severity failure;
	assert RAM(27090) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27090))))  severity failure;
	assert RAM(27091) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(27091))))  severity failure;
	assert RAM(27092) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(27092))))  severity failure;
	assert RAM(27093) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(27093))))  severity failure;
	assert RAM(27094) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27094))))  severity failure;
	assert RAM(27095) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27095))))  severity failure;
	assert RAM(27096) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27096))))  severity failure;
	assert RAM(27097) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(27097))))  severity failure;
	assert RAM(27098) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(27098))))  severity failure;
	assert RAM(27099) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(27099))))  severity failure;
	assert RAM(27100) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27100))))  severity failure;
	assert RAM(27101) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(27101))))  severity failure;
	assert RAM(27102) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27102))))  severity failure;
	assert RAM(27103) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(27103))))  severity failure;
	assert RAM(27104) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(27104))))  severity failure;
	assert RAM(27105) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(27105))))  severity failure;
	assert RAM(27106) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(27106))))  severity failure;
	assert RAM(27107) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(27107))))  severity failure;
	assert RAM(27108) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(27108))))  severity failure;
	assert RAM(27109) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27109))))  severity failure;
	assert RAM(27110) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27110))))  severity failure;
	assert RAM(27111) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(27111))))  severity failure;
	assert RAM(27112) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27112))))  severity failure;
	assert RAM(27113) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27113))))  severity failure;
	assert RAM(27114) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(27114))))  severity failure;
	assert RAM(27115) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(27115))))  severity failure;
	assert RAM(27116) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27116))))  severity failure;
	assert RAM(27117) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27117))))  severity failure;
	assert RAM(27118) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(27118))))  severity failure;
	assert RAM(27119) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27119))))  severity failure;
	assert RAM(27120) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(27120))))  severity failure;
	assert RAM(27121) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(27121))))  severity failure;
	assert RAM(27122) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27122))))  severity failure;
	assert RAM(27123) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(27123))))  severity failure;
	assert RAM(27124) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27124))))  severity failure;
	assert RAM(27125) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(27125))))  severity failure;
	assert RAM(27126) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(27126))))  severity failure;
	assert RAM(27127) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(27127))))  severity failure;
	assert RAM(27128) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(27128))))  severity failure;
	assert RAM(27129) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27129))))  severity failure;
	assert RAM(27130) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(27130))))  severity failure;
	assert RAM(27131) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(27131))))  severity failure;
	assert RAM(27132) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(27132))))  severity failure;
	assert RAM(27133) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(27133))))  severity failure;
	assert RAM(27134) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(27134))))  severity failure;
	assert RAM(27135) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27135))))  severity failure;
	assert RAM(27136) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(27136))))  severity failure;
	assert RAM(27137) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27137))))  severity failure;
	assert RAM(27138) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(27138))))  severity failure;
	assert RAM(27139) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(27139))))  severity failure;
	assert RAM(27140) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27140))))  severity failure;
	assert RAM(27141) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(27141))))  severity failure;
	assert RAM(27142) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27142))))  severity failure;
	assert RAM(27143) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27143))))  severity failure;
	assert RAM(27144) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(27144))))  severity failure;
	assert RAM(27145) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27145))))  severity failure;
	assert RAM(27146) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27146))))  severity failure;
	assert RAM(27147) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(27147))))  severity failure;
	assert RAM(27148) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(27148))))  severity failure;
	assert RAM(27149) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27149))))  severity failure;
	assert RAM(27150) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(27150))))  severity failure;
	assert RAM(27151) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(27151))))  severity failure;
	assert RAM(27152) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27152))))  severity failure;
	assert RAM(27153) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(27153))))  severity failure;
	assert RAM(27154) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(27154))))  severity failure;
	assert RAM(27155) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(27155))))  severity failure;
	assert RAM(27156) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(27156))))  severity failure;
	assert RAM(27157) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(27157))))  severity failure;
	assert RAM(27158) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(27158))))  severity failure;
	assert RAM(27159) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(27159))))  severity failure;
	assert RAM(27160) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(27160))))  severity failure;
	assert RAM(27161) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(27161))))  severity failure;
	assert RAM(27162) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27162))))  severity failure;
	assert RAM(27163) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27163))))  severity failure;
	assert RAM(27164) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(27164))))  severity failure;
	assert RAM(27165) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(27165))))  severity failure;
	assert RAM(27166) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(27166))))  severity failure;
	assert RAM(27167) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(27167))))  severity failure;
	assert RAM(27168) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(27168))))  severity failure;
	assert RAM(27169) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(27169))))  severity failure;
	assert RAM(27170) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(27170))))  severity failure;
	assert RAM(27171) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27171))))  severity failure;
	assert RAM(27172) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27172))))  severity failure;
	assert RAM(27173) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(27173))))  severity failure;
	assert RAM(27174) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27174))))  severity failure;
	assert RAM(27175) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(27175))))  severity failure;
	assert RAM(27176) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27176))))  severity failure;
	assert RAM(27177) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27177))))  severity failure;
	assert RAM(27178) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27178))))  severity failure;
	assert RAM(27179) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27179))))  severity failure;
	assert RAM(27180) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27180))))  severity failure;
	assert RAM(27181) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(27181))))  severity failure;
	assert RAM(27182) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(27182))))  severity failure;
	assert RAM(27183) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27183))))  severity failure;
	assert RAM(27184) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27184))))  severity failure;
	assert RAM(27185) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(27185))))  severity failure;
	assert RAM(27186) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(27186))))  severity failure;
	assert RAM(27187) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(27187))))  severity failure;
	assert RAM(27188) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27188))))  severity failure;
	assert RAM(27189) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27189))))  severity failure;
	assert RAM(27190) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(27190))))  severity failure;
	assert RAM(27191) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(27191))))  severity failure;
	assert RAM(27192) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(27192))))  severity failure;
	assert RAM(27193) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(27193))))  severity failure;
	assert RAM(27194) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(27194))))  severity failure;
	assert RAM(27195) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(27195))))  severity failure;
	assert RAM(27196) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27196))))  severity failure;
	assert RAM(27197) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(27197))))  severity failure;
	assert RAM(27198) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(27198))))  severity failure;
	assert RAM(27199) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(27199))))  severity failure;
	assert RAM(27200) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27200))))  severity failure;
	assert RAM(27201) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(27201))))  severity failure;
	assert RAM(27202) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(27202))))  severity failure;
	assert RAM(27203) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(27203))))  severity failure;
	assert RAM(27204) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27204))))  severity failure;
	assert RAM(27205) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(27205))))  severity failure;
	assert RAM(27206) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(27206))))  severity failure;
	assert RAM(27207) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(27207))))  severity failure;
	assert RAM(27208) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27208))))  severity failure;
	assert RAM(27209) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(27209))))  severity failure;
	assert RAM(27210) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(27210))))  severity failure;
	assert RAM(27211) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27211))))  severity failure;
	assert RAM(27212) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27212))))  severity failure;
	assert RAM(27213) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(27213))))  severity failure;
	assert RAM(27214) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(27214))))  severity failure;
	assert RAM(27215) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(27215))))  severity failure;
	assert RAM(27216) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(27216))))  severity failure;
	assert RAM(27217) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(27217))))  severity failure;
	assert RAM(27218) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(27218))))  severity failure;
	assert RAM(27219) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(27219))))  severity failure;
	assert RAM(27220) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27220))))  severity failure;
	assert RAM(27221) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(27221))))  severity failure;
	assert RAM(27222) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27222))))  severity failure;
	assert RAM(27223) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(27223))))  severity failure;
	assert RAM(27224) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27224))))  severity failure;
	assert RAM(27225) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(27225))))  severity failure;
	assert RAM(27226) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(27226))))  severity failure;
	assert RAM(27227) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27227))))  severity failure;
	assert RAM(27228) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(27228))))  severity failure;
	assert RAM(27229) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(27229))))  severity failure;
	assert RAM(27230) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(27230))))  severity failure;
	assert RAM(27231) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(27231))))  severity failure;
	assert RAM(27232) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27232))))  severity failure;
	assert RAM(27233) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(27233))))  severity failure;
	assert RAM(27234) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(27234))))  severity failure;
	assert RAM(27235) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(27235))))  severity failure;
	assert RAM(27236) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(27236))))  severity failure;
	assert RAM(27237) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(27237))))  severity failure;
	assert RAM(27238) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27238))))  severity failure;
	assert RAM(27239) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(27239))))  severity failure;
	assert RAM(27240) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(27240))))  severity failure;
	assert RAM(27241) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(27241))))  severity failure;
	assert RAM(27242) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27242))))  severity failure;
	assert RAM(27243) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27243))))  severity failure;
	assert RAM(27244) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(27244))))  severity failure;
	assert RAM(27245) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(27245))))  severity failure;
	assert RAM(27246) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(27246))))  severity failure;
	assert RAM(27247) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(27247))))  severity failure;
	assert RAM(27248) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(27248))))  severity failure;
	assert RAM(27249) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(27249))))  severity failure;
	assert RAM(27250) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(27250))))  severity failure;
	assert RAM(27251) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27251))))  severity failure;
	assert RAM(27252) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(27252))))  severity failure;
	assert RAM(27253) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(27253))))  severity failure;
	assert RAM(27254) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(27254))))  severity failure;
	assert RAM(27255) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(27255))))  severity failure;
	assert RAM(27256) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(27256))))  severity failure;
	assert RAM(27257) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(27257))))  severity failure;
	assert RAM(27258) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(27258))))  severity failure;
	assert RAM(27259) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(27259))))  severity failure;
	assert RAM(27260) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27260))))  severity failure;
	assert RAM(27261) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27261))))  severity failure;
	assert RAM(27262) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(27262))))  severity failure;
	assert RAM(27263) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(27263))))  severity failure;
	assert RAM(27264) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27264))))  severity failure;
	assert RAM(27265) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(27265))))  severity failure;
	assert RAM(27266) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27266))))  severity failure;
	assert RAM(27267) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(27267))))  severity failure;
	assert RAM(27268) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(27268))))  severity failure;
	assert RAM(27269) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27269))))  severity failure;
	assert RAM(27270) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(27270))))  severity failure;
	assert RAM(27271) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(27271))))  severity failure;
	assert RAM(27272) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27272))))  severity failure;
	assert RAM(27273) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(27273))))  severity failure;
	assert RAM(27274) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(27274))))  severity failure;
	assert RAM(27275) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27275))))  severity failure;
	assert RAM(27276) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27276))))  severity failure;
	assert RAM(27277) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(27277))))  severity failure;
	assert RAM(27278) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(27278))))  severity failure;
	assert RAM(27279) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27279))))  severity failure;
	assert RAM(27280) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(27280))))  severity failure;
	assert RAM(27281) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(27281))))  severity failure;
	assert RAM(27282) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(27282))))  severity failure;
	assert RAM(27283) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27283))))  severity failure;
	assert RAM(27284) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(27284))))  severity failure;
	assert RAM(27285) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(27285))))  severity failure;
	assert RAM(27286) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(27286))))  severity failure;
	assert RAM(27287) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(27287))))  severity failure;
	assert RAM(27288) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(27288))))  severity failure;
	assert RAM(27289) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(27289))))  severity failure;
	assert RAM(27290) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(27290))))  severity failure;
	assert RAM(27291) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(27291))))  severity failure;
	assert RAM(27292) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(27292))))  severity failure;
	assert RAM(27293) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(27293))))  severity failure;
	assert RAM(27294) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(27294))))  severity failure;
	assert RAM(27295) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(27295))))  severity failure;
	assert RAM(27296) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(27296))))  severity failure;
	assert RAM(27297) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27297))))  severity failure;
	assert RAM(27298) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27298))))  severity failure;
	assert RAM(27299) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(27299))))  severity failure;
	assert RAM(27300) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27300))))  severity failure;
	assert RAM(27301) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27301))))  severity failure;
	assert RAM(27302) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(27302))))  severity failure;
	assert RAM(27303) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27303))))  severity failure;
	assert RAM(27304) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(27304))))  severity failure;
	assert RAM(27305) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27305))))  severity failure;
	assert RAM(27306) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(27306))))  severity failure;
	assert RAM(27307) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27307))))  severity failure;
	assert RAM(27308) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(27308))))  severity failure;
	assert RAM(27309) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(27309))))  severity failure;
	assert RAM(27310) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27310))))  severity failure;
	assert RAM(27311) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(27311))))  severity failure;
	assert RAM(27312) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27312))))  severity failure;
	assert RAM(27313) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(27313))))  severity failure;
	assert RAM(27314) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(27314))))  severity failure;
	assert RAM(27315) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(27315))))  severity failure;
	assert RAM(27316) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(27316))))  severity failure;
	assert RAM(27317) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27317))))  severity failure;
	assert RAM(27318) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27318))))  severity failure;
	assert RAM(27319) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(27319))))  severity failure;
	assert RAM(27320) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27320))))  severity failure;
	assert RAM(27321) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27321))))  severity failure;
	assert RAM(27322) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27322))))  severity failure;
	assert RAM(27323) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(27323))))  severity failure;
	assert RAM(27324) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(27324))))  severity failure;
	assert RAM(27325) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(27325))))  severity failure;
	assert RAM(27326) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27326))))  severity failure;
	assert RAM(27327) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(27327))))  severity failure;
	assert RAM(27328) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(27328))))  severity failure;
	assert RAM(27329) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27329))))  severity failure;
	assert RAM(27330) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(27330))))  severity failure;
	assert RAM(27331) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27331))))  severity failure;
	assert RAM(27332) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(27332))))  severity failure;
	assert RAM(27333) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(27333))))  severity failure;
	assert RAM(27334) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(27334))))  severity failure;
	assert RAM(27335) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27335))))  severity failure;
	assert RAM(27336) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27336))))  severity failure;
	assert RAM(27337) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27337))))  severity failure;
	assert RAM(27338) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(27338))))  severity failure;
	assert RAM(27339) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27339))))  severity failure;
	assert RAM(27340) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(27340))))  severity failure;
	assert RAM(27341) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27341))))  severity failure;
	assert RAM(27342) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(27342))))  severity failure;
	assert RAM(27343) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(27343))))  severity failure;
	assert RAM(27344) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(27344))))  severity failure;
	assert RAM(27345) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27345))))  severity failure;
	assert RAM(27346) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(27346))))  severity failure;
	assert RAM(27347) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27347))))  severity failure;
	assert RAM(27348) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27348))))  severity failure;
	assert RAM(27349) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(27349))))  severity failure;
	assert RAM(27350) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27350))))  severity failure;
	assert RAM(27351) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(27351))))  severity failure;
	assert RAM(27352) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(27352))))  severity failure;
	assert RAM(27353) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(27353))))  severity failure;
	assert RAM(27354) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(27354))))  severity failure;
	assert RAM(27355) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(27355))))  severity failure;
	assert RAM(27356) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(27356))))  severity failure;
	assert RAM(27357) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27357))))  severity failure;
	assert RAM(27358) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27358))))  severity failure;
	assert RAM(27359) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(27359))))  severity failure;
	assert RAM(27360) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27360))))  severity failure;
	assert RAM(27361) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(27361))))  severity failure;
	assert RAM(27362) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(27362))))  severity failure;
	assert RAM(27363) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(27363))))  severity failure;
	assert RAM(27364) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(27364))))  severity failure;
	assert RAM(27365) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(27365))))  severity failure;
	assert RAM(27366) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(27366))))  severity failure;
	assert RAM(27367) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(27367))))  severity failure;
	assert RAM(27368) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27368))))  severity failure;
	assert RAM(27369) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(27369))))  severity failure;
	assert RAM(27370) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(27370))))  severity failure;
	assert RAM(27371) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(27371))))  severity failure;
	assert RAM(27372) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27372))))  severity failure;
	assert RAM(27373) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27373))))  severity failure;
	assert RAM(27374) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27374))))  severity failure;
	assert RAM(27375) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27375))))  severity failure;
	assert RAM(27376) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27376))))  severity failure;
	assert RAM(27377) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27377))))  severity failure;
	assert RAM(27378) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(27378))))  severity failure;
	assert RAM(27379) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27379))))  severity failure;
	assert RAM(27380) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27380))))  severity failure;
	assert RAM(27381) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27381))))  severity failure;
	assert RAM(27382) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27382))))  severity failure;
	assert RAM(27383) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(27383))))  severity failure;
	assert RAM(27384) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(27384))))  severity failure;
	assert RAM(27385) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(27385))))  severity failure;
	assert RAM(27386) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27386))))  severity failure;
	assert RAM(27387) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27387))))  severity failure;
	assert RAM(27388) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27388))))  severity failure;
	assert RAM(27389) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27389))))  severity failure;
	assert RAM(27390) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(27390))))  severity failure;
	assert RAM(27391) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(27391))))  severity failure;
	assert RAM(27392) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(27392))))  severity failure;
	assert RAM(27393) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(27393))))  severity failure;
	assert RAM(27394) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(27394))))  severity failure;
	assert RAM(27395) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27395))))  severity failure;
	assert RAM(27396) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27396))))  severity failure;
	assert RAM(27397) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(27397))))  severity failure;
	assert RAM(27398) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(27398))))  severity failure;
	assert RAM(27399) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27399))))  severity failure;
	assert RAM(27400) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(27400))))  severity failure;
	assert RAM(27401) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27401))))  severity failure;
	assert RAM(27402) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(27402))))  severity failure;
	assert RAM(27403) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(27403))))  severity failure;
	assert RAM(27404) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27404))))  severity failure;
	assert RAM(27405) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27405))))  severity failure;
	assert RAM(27406) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(27406))))  severity failure;
	assert RAM(27407) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(27407))))  severity failure;
	assert RAM(27408) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(27408))))  severity failure;
	assert RAM(27409) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(27409))))  severity failure;
	assert RAM(27410) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(27410))))  severity failure;
	assert RAM(27411) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(27411))))  severity failure;
	assert RAM(27412) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27412))))  severity failure;
	assert RAM(27413) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(27413))))  severity failure;
	assert RAM(27414) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(27414))))  severity failure;
	assert RAM(27415) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(27415))))  severity failure;
	assert RAM(27416) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27416))))  severity failure;
	assert RAM(27417) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27417))))  severity failure;
	assert RAM(27418) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(27418))))  severity failure;
	assert RAM(27419) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(27419))))  severity failure;
	assert RAM(27420) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(27420))))  severity failure;
	assert RAM(27421) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27421))))  severity failure;
	assert RAM(27422) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27422))))  severity failure;
	assert RAM(27423) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(27423))))  severity failure;
	assert RAM(27424) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(27424))))  severity failure;
	assert RAM(27425) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27425))))  severity failure;
	assert RAM(27426) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(27426))))  severity failure;
	assert RAM(27427) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(27427))))  severity failure;
	assert RAM(27428) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(27428))))  severity failure;
	assert RAM(27429) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(27429))))  severity failure;
	assert RAM(27430) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(27430))))  severity failure;
	assert RAM(27431) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(27431))))  severity failure;
	assert RAM(27432) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(27432))))  severity failure;
	assert RAM(27433) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(27433))))  severity failure;
	assert RAM(27434) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(27434))))  severity failure;
	assert RAM(27435) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(27435))))  severity failure;
	assert RAM(27436) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(27436))))  severity failure;
	assert RAM(27437) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(27437))))  severity failure;
	assert RAM(27438) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27438))))  severity failure;
	assert RAM(27439) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(27439))))  severity failure;
	assert RAM(27440) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(27440))))  severity failure;
	assert RAM(27441) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27441))))  severity failure;
	assert RAM(27442) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(27442))))  severity failure;
	assert RAM(27443) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(27443))))  severity failure;
	assert RAM(27444) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(27444))))  severity failure;
	assert RAM(27445) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(27445))))  severity failure;
	assert RAM(27446) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(27446))))  severity failure;
	assert RAM(27447) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(27447))))  severity failure;
	assert RAM(27448) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27448))))  severity failure;
	assert RAM(27449) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(27449))))  severity failure;
	assert RAM(27450) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(27450))))  severity failure;
	assert RAM(27451) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(27451))))  severity failure;
	assert RAM(27452) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(27452))))  severity failure;
	assert RAM(27453) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(27453))))  severity failure;
	assert RAM(27454) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(27454))))  severity failure;
	assert RAM(27455) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(27455))))  severity failure;
	assert RAM(27456) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(27456))))  severity failure;
	assert RAM(27457) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(27457))))  severity failure;
	assert RAM(27458) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27458))))  severity failure;
	assert RAM(27459) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(27459))))  severity failure;
	assert RAM(27460) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(27460))))  severity failure;
	assert RAM(27461) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(27461))))  severity failure;
	assert RAM(27462) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27462))))  severity failure;
	assert RAM(27463) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27463))))  severity failure;
	assert RAM(27464) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27464))))  severity failure;
	assert RAM(27465) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27465))))  severity failure;
	assert RAM(27466) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27466))))  severity failure;
	assert RAM(27467) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(27467))))  severity failure;
	assert RAM(27468) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(27468))))  severity failure;
	assert RAM(27469) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(27469))))  severity failure;
	assert RAM(27470) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(27470))))  severity failure;
	assert RAM(27471) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27471))))  severity failure;
	assert RAM(27472) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(27472))))  severity failure;
	assert RAM(27473) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27473))))  severity failure;
	assert RAM(27474) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27474))))  severity failure;
	assert RAM(27475) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(27475))))  severity failure;
	assert RAM(27476) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(27476))))  severity failure;
	assert RAM(27477) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(27477))))  severity failure;
	assert RAM(27478) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(27478))))  severity failure;
	assert RAM(27479) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27479))))  severity failure;
	assert RAM(27480) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(27480))))  severity failure;
	assert RAM(27481) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(27481))))  severity failure;
	assert RAM(27482) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(27482))))  severity failure;
	assert RAM(27483) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(27483))))  severity failure;
	assert RAM(27484) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27484))))  severity failure;
	assert RAM(27485) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(27485))))  severity failure;
	assert RAM(27486) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27486))))  severity failure;
	assert RAM(27487) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27487))))  severity failure;
	assert RAM(27488) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27488))))  severity failure;
	assert RAM(27489) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(27489))))  severity failure;
	assert RAM(27490) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(27490))))  severity failure;
	assert RAM(27491) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(27491))))  severity failure;
	assert RAM(27492) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(27492))))  severity failure;
	assert RAM(27493) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(27493))))  severity failure;
	assert RAM(27494) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27494))))  severity failure;
	assert RAM(27495) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(27495))))  severity failure;
	assert RAM(27496) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27496))))  severity failure;
	assert RAM(27497) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(27497))))  severity failure;
	assert RAM(27498) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(27498))))  severity failure;
	assert RAM(27499) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(27499))))  severity failure;
	assert RAM(27500) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(27500))))  severity failure;
	assert RAM(27501) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27501))))  severity failure;
	assert RAM(27502) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(27502))))  severity failure;
	assert RAM(27503) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(27503))))  severity failure;
	assert RAM(27504) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27504))))  severity failure;
	assert RAM(27505) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27505))))  severity failure;
	assert RAM(27506) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(27506))))  severity failure;
	assert RAM(27507) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(27507))))  severity failure;
	assert RAM(27508) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(27508))))  severity failure;
	assert RAM(27509) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27509))))  severity failure;
	assert RAM(27510) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27510))))  severity failure;
	assert RAM(27511) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(27511))))  severity failure;
	assert RAM(27512) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27512))))  severity failure;
	assert RAM(27513) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(27513))))  severity failure;
	assert RAM(27514) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(27514))))  severity failure;
	assert RAM(27515) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27515))))  severity failure;
	assert RAM(27516) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27516))))  severity failure;
	assert RAM(27517) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(27517))))  severity failure;
	assert RAM(27518) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27518))))  severity failure;
	assert RAM(27519) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27519))))  severity failure;
	assert RAM(27520) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27520))))  severity failure;
	assert RAM(27521) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27521))))  severity failure;
	assert RAM(27522) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(27522))))  severity failure;
	assert RAM(27523) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27523))))  severity failure;
	assert RAM(27524) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(27524))))  severity failure;
	assert RAM(27525) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(27525))))  severity failure;
	assert RAM(27526) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(27526))))  severity failure;
	assert RAM(27527) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(27527))))  severity failure;
	assert RAM(27528) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(27528))))  severity failure;
	assert RAM(27529) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(27529))))  severity failure;
	assert RAM(27530) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27530))))  severity failure;
	assert RAM(27531) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(27531))))  severity failure;
	assert RAM(27532) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(27532))))  severity failure;
	assert RAM(27533) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(27533))))  severity failure;
	assert RAM(27534) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(27534))))  severity failure;
	assert RAM(27535) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(27535))))  severity failure;
	assert RAM(27536) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27536))))  severity failure;
	assert RAM(27537) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(27537))))  severity failure;
	assert RAM(27538) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27538))))  severity failure;
	assert RAM(27539) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(27539))))  severity failure;
	assert RAM(27540) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(27540))))  severity failure;
	assert RAM(27541) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27541))))  severity failure;
	assert RAM(27542) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27542))))  severity failure;
	assert RAM(27543) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(27543))))  severity failure;
	assert RAM(27544) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(27544))))  severity failure;
	assert RAM(27545) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27545))))  severity failure;
	assert RAM(27546) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(27546))))  severity failure;
	assert RAM(27547) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(27547))))  severity failure;
	assert RAM(27548) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(27548))))  severity failure;
	assert RAM(27549) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27549))))  severity failure;
	assert RAM(27550) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27550))))  severity failure;
	assert RAM(27551) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(27551))))  severity failure;
	assert RAM(27552) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(27552))))  severity failure;
	assert RAM(27553) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(27553))))  severity failure;
	assert RAM(27554) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27554))))  severity failure;
	assert RAM(27555) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(27555))))  severity failure;
	assert RAM(27556) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27556))))  severity failure;
	assert RAM(27557) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(27557))))  severity failure;
	assert RAM(27558) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(27558))))  severity failure;
	assert RAM(27559) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(27559))))  severity failure;
	assert RAM(27560) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(27560))))  severity failure;
	assert RAM(27561) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(27561))))  severity failure;
	assert RAM(27562) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(27562))))  severity failure;
	assert RAM(27563) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27563))))  severity failure;
	assert RAM(27564) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(27564))))  severity failure;
	assert RAM(27565) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27565))))  severity failure;
	assert RAM(27566) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27566))))  severity failure;
	assert RAM(27567) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(27567))))  severity failure;
	assert RAM(27568) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(27568))))  severity failure;
	assert RAM(27569) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27569))))  severity failure;
	assert RAM(27570) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(27570))))  severity failure;
	assert RAM(27571) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27571))))  severity failure;
	assert RAM(27572) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27572))))  severity failure;
	assert RAM(27573) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27573))))  severity failure;
	assert RAM(27574) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27574))))  severity failure;
	assert RAM(27575) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27575))))  severity failure;
	assert RAM(27576) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27576))))  severity failure;
	assert RAM(27577) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(27577))))  severity failure;
	assert RAM(27578) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(27578))))  severity failure;
	assert RAM(27579) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(27579))))  severity failure;
	assert RAM(27580) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(27580))))  severity failure;
	assert RAM(27581) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(27581))))  severity failure;
	assert RAM(27582) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(27582))))  severity failure;
	assert RAM(27583) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(27583))))  severity failure;
	assert RAM(27584) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27584))))  severity failure;
	assert RAM(27585) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(27585))))  severity failure;
	assert RAM(27586) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(27586))))  severity failure;
	assert RAM(27587) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(27587))))  severity failure;
	assert RAM(27588) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27588))))  severity failure;
	assert RAM(27589) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27589))))  severity failure;
	assert RAM(27590) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(27590))))  severity failure;
	assert RAM(27591) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(27591))))  severity failure;
	assert RAM(27592) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27592))))  severity failure;
	assert RAM(27593) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(27593))))  severity failure;
	assert RAM(27594) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(27594))))  severity failure;
	assert RAM(27595) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(27595))))  severity failure;
	assert RAM(27596) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27596))))  severity failure;
	assert RAM(27597) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(27597))))  severity failure;
	assert RAM(27598) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27598))))  severity failure;
	assert RAM(27599) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(27599))))  severity failure;
	assert RAM(27600) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27600))))  severity failure;
	assert RAM(27601) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(27601))))  severity failure;
	assert RAM(27602) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27602))))  severity failure;
	assert RAM(27603) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(27603))))  severity failure;
	assert RAM(27604) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(27604))))  severity failure;
	assert RAM(27605) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(27605))))  severity failure;
	assert RAM(27606) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(27606))))  severity failure;
	assert RAM(27607) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27607))))  severity failure;
	assert RAM(27608) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(27608))))  severity failure;
	assert RAM(27609) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27609))))  severity failure;
	assert RAM(27610) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(27610))))  severity failure;
	assert RAM(27611) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27611))))  severity failure;
	assert RAM(27612) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(27612))))  severity failure;
	assert RAM(27613) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(27613))))  severity failure;
	assert RAM(27614) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(27614))))  severity failure;
	assert RAM(27615) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27615))))  severity failure;
	assert RAM(27616) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(27616))))  severity failure;
	assert RAM(27617) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(27617))))  severity failure;
	assert RAM(27618) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(27618))))  severity failure;
	assert RAM(27619) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(27619))))  severity failure;
	assert RAM(27620) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27620))))  severity failure;
	assert RAM(27621) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(27621))))  severity failure;
	assert RAM(27622) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(27622))))  severity failure;
	assert RAM(27623) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(27623))))  severity failure;
	assert RAM(27624) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(27624))))  severity failure;
	assert RAM(27625) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(27625))))  severity failure;
	assert RAM(27626) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(27626))))  severity failure;
	assert RAM(27627) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(27627))))  severity failure;
	assert RAM(27628) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(27628))))  severity failure;
	assert RAM(27629) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(27629))))  severity failure;
	assert RAM(27630) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27630))))  severity failure;
	assert RAM(27631) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(27631))))  severity failure;
	assert RAM(27632) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27632))))  severity failure;
	assert RAM(27633) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(27633))))  severity failure;
	assert RAM(27634) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(27634))))  severity failure;
	assert RAM(27635) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(27635))))  severity failure;
	assert RAM(27636) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(27636))))  severity failure;
	assert RAM(27637) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(27637))))  severity failure;
	assert RAM(27638) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27638))))  severity failure;
	assert RAM(27639) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(27639))))  severity failure;
	assert RAM(27640) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(27640))))  severity failure;
	assert RAM(27641) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27641))))  severity failure;
	assert RAM(27642) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(27642))))  severity failure;
	assert RAM(27643) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(27643))))  severity failure;
	assert RAM(27644) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(27644))))  severity failure;
	assert RAM(27645) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27645))))  severity failure;
	assert RAM(27646) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(27646))))  severity failure;
	assert RAM(27647) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(27647))))  severity failure;
	assert RAM(27648) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(27648))))  severity failure;
	assert RAM(27649) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(27649))))  severity failure;
	assert RAM(27650) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(27650))))  severity failure;
	assert RAM(27651) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(27651))))  severity failure;
	assert RAM(27652) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(27652))))  severity failure;
	assert RAM(27653) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27653))))  severity failure;
	assert RAM(27654) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(27654))))  severity failure;
	assert RAM(27655) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27655))))  severity failure;
	assert RAM(27656) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27656))))  severity failure;
	assert RAM(27657) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27657))))  severity failure;
	assert RAM(27658) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(27658))))  severity failure;
	assert RAM(27659) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(27659))))  severity failure;
	assert RAM(27660) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(27660))))  severity failure;
	assert RAM(27661) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(27661))))  severity failure;
	assert RAM(27662) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27662))))  severity failure;
	assert RAM(27663) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27663))))  severity failure;
	assert RAM(27664) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(27664))))  severity failure;
	assert RAM(27665) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27665))))  severity failure;
	assert RAM(27666) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27666))))  severity failure;
	assert RAM(27667) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(27667))))  severity failure;
	assert RAM(27668) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(27668))))  severity failure;
	assert RAM(27669) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(27669))))  severity failure;
	assert RAM(27670) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(27670))))  severity failure;
	assert RAM(27671) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27671))))  severity failure;
	assert RAM(27672) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27672))))  severity failure;
	assert RAM(27673) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(27673))))  severity failure;
	assert RAM(27674) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(27674))))  severity failure;
	assert RAM(27675) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(27675))))  severity failure;
	assert RAM(27676) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27676))))  severity failure;
	assert RAM(27677) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(27677))))  severity failure;
	assert RAM(27678) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(27678))))  severity failure;
	assert RAM(27679) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(27679))))  severity failure;
	assert RAM(27680) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(27680))))  severity failure;
	assert RAM(27681) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(27681))))  severity failure;
	assert RAM(27682) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(27682))))  severity failure;
	assert RAM(27683) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27683))))  severity failure;
	assert RAM(27684) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(27684))))  severity failure;
	assert RAM(27685) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27685))))  severity failure;
	assert RAM(27686) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(27686))))  severity failure;
	assert RAM(27687) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27687))))  severity failure;
	assert RAM(27688) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(27688))))  severity failure;
	assert RAM(27689) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27689))))  severity failure;
	assert RAM(27690) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(27690))))  severity failure;
	assert RAM(27691) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(27691))))  severity failure;
	assert RAM(27692) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(27692))))  severity failure;
	assert RAM(27693) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27693))))  severity failure;
	assert RAM(27694) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(27694))))  severity failure;
	assert RAM(27695) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(27695))))  severity failure;
	assert RAM(27696) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27696))))  severity failure;
	assert RAM(27697) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(27697))))  severity failure;
	assert RAM(27698) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(27698))))  severity failure;
	assert RAM(27699) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(27699))))  severity failure;
	assert RAM(27700) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(27700))))  severity failure;
	assert RAM(27701) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(27701))))  severity failure;
	assert RAM(27702) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27702))))  severity failure;
	assert RAM(27703) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(27703))))  severity failure;
	assert RAM(27704) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27704))))  severity failure;
	assert RAM(27705) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(27705))))  severity failure;
	assert RAM(27706) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27706))))  severity failure;
	assert RAM(27707) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(27707))))  severity failure;
	assert RAM(27708) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(27708))))  severity failure;
	assert RAM(27709) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(27709))))  severity failure;
	assert RAM(27710) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(27710))))  severity failure;
	assert RAM(27711) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(27711))))  severity failure;
	assert RAM(27712) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(27712))))  severity failure;
	assert RAM(27713) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(27713))))  severity failure;
	assert RAM(27714) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(27714))))  severity failure;
	assert RAM(27715) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27715))))  severity failure;
	assert RAM(27716) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(27716))))  severity failure;
	assert RAM(27717) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(27717))))  severity failure;
	assert RAM(27718) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27718))))  severity failure;
	assert RAM(27719) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(27719))))  severity failure;
	assert RAM(27720) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(27720))))  severity failure;
	assert RAM(27721) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27721))))  severity failure;
	assert RAM(27722) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(27722))))  severity failure;
	assert RAM(27723) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(27723))))  severity failure;
	assert RAM(27724) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(27724))))  severity failure;
	assert RAM(27725) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(27725))))  severity failure;
	assert RAM(27726) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27726))))  severity failure;
	assert RAM(27727) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(27727))))  severity failure;
	assert RAM(27728) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(27728))))  severity failure;
	assert RAM(27729) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27729))))  severity failure;
	assert RAM(27730) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(27730))))  severity failure;
	assert RAM(27731) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(27731))))  severity failure;
	assert RAM(27732) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27732))))  severity failure;
	assert RAM(27733) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27733))))  severity failure;
	assert RAM(27734) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(27734))))  severity failure;
	assert RAM(27735) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(27735))))  severity failure;
	assert RAM(27736) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(27736))))  severity failure;
	assert RAM(27737) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(27737))))  severity failure;
	assert RAM(27738) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(27738))))  severity failure;
	assert RAM(27739) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(27739))))  severity failure;
	assert RAM(27740) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(27740))))  severity failure;
	assert RAM(27741) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27741))))  severity failure;
	assert RAM(27742) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(27742))))  severity failure;
	assert RAM(27743) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27743))))  severity failure;
	assert RAM(27744) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(27744))))  severity failure;
	assert RAM(27745) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27745))))  severity failure;
	assert RAM(27746) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(27746))))  severity failure;
	assert RAM(27747) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27747))))  severity failure;
	assert RAM(27748) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(27748))))  severity failure;
	assert RAM(27749) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(27749))))  severity failure;
	assert RAM(27750) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(27750))))  severity failure;
	assert RAM(27751) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(27751))))  severity failure;
	assert RAM(27752) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27752))))  severity failure;
	assert RAM(27753) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(27753))))  severity failure;
	assert RAM(27754) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(27754))))  severity failure;
	assert RAM(27755) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27755))))  severity failure;
	assert RAM(27756) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(27756))))  severity failure;
	assert RAM(27757) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(27757))))  severity failure;
	assert RAM(27758) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(27758))))  severity failure;
	assert RAM(27759) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(27759))))  severity failure;
	assert RAM(27760) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(27760))))  severity failure;
	assert RAM(27761) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(27761))))  severity failure;
	assert RAM(27762) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27762))))  severity failure;
	assert RAM(27763) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(27763))))  severity failure;
	assert RAM(27764) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(27764))))  severity failure;
	assert RAM(27765) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(27765))))  severity failure;
	assert RAM(27766) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(27766))))  severity failure;
	assert RAM(27767) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27767))))  severity failure;
	assert RAM(27768) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(27768))))  severity failure;
	assert RAM(27769) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27769))))  severity failure;
	assert RAM(27770) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(27770))))  severity failure;
	assert RAM(27771) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(27771))))  severity failure;
	assert RAM(27772) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(27772))))  severity failure;
	assert RAM(27773) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(27773))))  severity failure;
	assert RAM(27774) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(27774))))  severity failure;
	assert RAM(27775) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(27775))))  severity failure;
	assert RAM(27776) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(27776))))  severity failure;
	assert RAM(27777) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27777))))  severity failure;
	assert RAM(27778) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(27778))))  severity failure;
	assert RAM(27779) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(27779))))  severity failure;
	assert RAM(27780) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(27780))))  severity failure;
	assert RAM(27781) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(27781))))  severity failure;
	assert RAM(27782) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(27782))))  severity failure;
	assert RAM(27783) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27783))))  severity failure;
	assert RAM(27784) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27784))))  severity failure;
	assert RAM(27785) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(27785))))  severity failure;
	assert RAM(27786) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(27786))))  severity failure;
	assert RAM(27787) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(27787))))  severity failure;
	assert RAM(27788) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(27788))))  severity failure;
	assert RAM(27789) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(27789))))  severity failure;
	assert RAM(27790) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(27790))))  severity failure;
	assert RAM(27791) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27791))))  severity failure;
	assert RAM(27792) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27792))))  severity failure;
	assert RAM(27793) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(27793))))  severity failure;
	assert RAM(27794) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(27794))))  severity failure;
	assert RAM(27795) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27795))))  severity failure;
	assert RAM(27796) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(27796))))  severity failure;
	assert RAM(27797) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(27797))))  severity failure;
	assert RAM(27798) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(27798))))  severity failure;
	assert RAM(27799) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27799))))  severity failure;
	assert RAM(27800) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(27800))))  severity failure;
	assert RAM(27801) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(27801))))  severity failure;
	assert RAM(27802) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(27802))))  severity failure;
	assert RAM(27803) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27803))))  severity failure;
	assert RAM(27804) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(27804))))  severity failure;
	assert RAM(27805) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(27805))))  severity failure;
	assert RAM(27806) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(27806))))  severity failure;
	assert RAM(27807) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27807))))  severity failure;
	assert RAM(27808) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27808))))  severity failure;
	assert RAM(27809) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(27809))))  severity failure;
	assert RAM(27810) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27810))))  severity failure;
	assert RAM(27811) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27811))))  severity failure;
	assert RAM(27812) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(27812))))  severity failure;
	assert RAM(27813) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(27813))))  severity failure;
	assert RAM(27814) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(27814))))  severity failure;
	assert RAM(27815) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27815))))  severity failure;
	assert RAM(27816) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(27816))))  severity failure;
	assert RAM(27817) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(27817))))  severity failure;
	assert RAM(27818) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27818))))  severity failure;
	assert RAM(27819) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(27819))))  severity failure;
	assert RAM(27820) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27820))))  severity failure;
	assert RAM(27821) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27821))))  severity failure;
	assert RAM(27822) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(27822))))  severity failure;
	assert RAM(27823) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(27823))))  severity failure;
	assert RAM(27824) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27824))))  severity failure;
	assert RAM(27825) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(27825))))  severity failure;
	assert RAM(27826) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27826))))  severity failure;
	assert RAM(27827) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(27827))))  severity failure;
	assert RAM(27828) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(27828))))  severity failure;
	assert RAM(27829) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27829))))  severity failure;
	assert RAM(27830) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(27830))))  severity failure;
	assert RAM(27831) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27831))))  severity failure;
	assert RAM(27832) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27832))))  severity failure;
	assert RAM(27833) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(27833))))  severity failure;
	assert RAM(27834) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27834))))  severity failure;
	assert RAM(27835) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(27835))))  severity failure;
	assert RAM(27836) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(27836))))  severity failure;
	assert RAM(27837) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(27837))))  severity failure;
	assert RAM(27838) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(27838))))  severity failure;
	assert RAM(27839) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(27839))))  severity failure;
	assert RAM(27840) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(27840))))  severity failure;
	assert RAM(27841) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(27841))))  severity failure;
	assert RAM(27842) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(27842))))  severity failure;
	assert RAM(27843) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(27843))))  severity failure;
	assert RAM(27844) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(27844))))  severity failure;
	assert RAM(27845) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(27845))))  severity failure;
	assert RAM(27846) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(27846))))  severity failure;
	assert RAM(27847) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(27847))))  severity failure;
	assert RAM(27848) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27848))))  severity failure;
	assert RAM(27849) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27849))))  severity failure;
	assert RAM(27850) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(27850))))  severity failure;
	assert RAM(27851) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(27851))))  severity failure;
	assert RAM(27852) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(27852))))  severity failure;
	assert RAM(27853) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(27853))))  severity failure;
	assert RAM(27854) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27854))))  severity failure;
	assert RAM(27855) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(27855))))  severity failure;
	assert RAM(27856) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27856))))  severity failure;
	assert RAM(27857) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(27857))))  severity failure;
	assert RAM(27858) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27858))))  severity failure;
	assert RAM(27859) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(27859))))  severity failure;
	assert RAM(27860) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(27860))))  severity failure;
	assert RAM(27861) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27861))))  severity failure;
	assert RAM(27862) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27862))))  severity failure;
	assert RAM(27863) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(27863))))  severity failure;
	assert RAM(27864) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(27864))))  severity failure;
	assert RAM(27865) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(27865))))  severity failure;
	assert RAM(27866) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(27866))))  severity failure;
	assert RAM(27867) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(27867))))  severity failure;
	assert RAM(27868) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(27868))))  severity failure;
	assert RAM(27869) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(27869))))  severity failure;
	assert RAM(27870) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(27870))))  severity failure;
	assert RAM(27871) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(27871))))  severity failure;
	assert RAM(27872) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(27872))))  severity failure;
	assert RAM(27873) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(27873))))  severity failure;
	assert RAM(27874) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(27874))))  severity failure;
	assert RAM(27875) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27875))))  severity failure;
	assert RAM(27876) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(27876))))  severity failure;
	assert RAM(27877) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(27877))))  severity failure;
	assert RAM(27878) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(27878))))  severity failure;
	assert RAM(27879) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(27879))))  severity failure;
	assert RAM(27880) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(27880))))  severity failure;
	assert RAM(27881) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(27881))))  severity failure;
	assert RAM(27882) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27882))))  severity failure;
	assert RAM(27883) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(27883))))  severity failure;
	assert RAM(27884) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27884))))  severity failure;
	assert RAM(27885) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(27885))))  severity failure;
	assert RAM(27886) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(27886))))  severity failure;
	assert RAM(27887) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(27887))))  severity failure;
	assert RAM(27888) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(27888))))  severity failure;
	assert RAM(27889) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(27889))))  severity failure;
	assert RAM(27890) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(27890))))  severity failure;
	assert RAM(27891) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(27891))))  severity failure;
	assert RAM(27892) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(27892))))  severity failure;
	assert RAM(27893) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(27893))))  severity failure;
	assert RAM(27894) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(27894))))  severity failure;
	assert RAM(27895) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(27895))))  severity failure;
	assert RAM(27896) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(27896))))  severity failure;
	assert RAM(27897) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(27897))))  severity failure;
	assert RAM(27898) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(27898))))  severity failure;
	assert RAM(27899) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(27899))))  severity failure;
	assert RAM(27900) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(27900))))  severity failure;
	assert RAM(27901) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(27901))))  severity failure;
	assert RAM(27902) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(27902))))  severity failure;
	assert RAM(27903) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(27903))))  severity failure;
	assert RAM(27904) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(27904))))  severity failure;
	assert RAM(27905) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27905))))  severity failure;
	assert RAM(27906) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27906))))  severity failure;
	assert RAM(27907) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27907))))  severity failure;
	assert RAM(27908) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(27908))))  severity failure;
	assert RAM(27909) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(27909))))  severity failure;
	assert RAM(27910) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(27910))))  severity failure;
	assert RAM(27911) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(27911))))  severity failure;
	assert RAM(27912) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(27912))))  severity failure;
	assert RAM(27913) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(27913))))  severity failure;
	assert RAM(27914) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(27914))))  severity failure;
	assert RAM(27915) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(27915))))  severity failure;
	assert RAM(27916) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(27916))))  severity failure;
	assert RAM(27917) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(27917))))  severity failure;
	assert RAM(27918) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(27918))))  severity failure;
	assert RAM(27919) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(27919))))  severity failure;
	assert RAM(27920) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(27920))))  severity failure;
	assert RAM(27921) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(27921))))  severity failure;
	assert RAM(27922) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(27922))))  severity failure;
	assert RAM(27923) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(27923))))  severity failure;
	assert RAM(27924) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(27924))))  severity failure;
	assert RAM(27925) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(27925))))  severity failure;
	assert RAM(27926) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(27926))))  severity failure;
	assert RAM(27927) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(27927))))  severity failure;
	assert RAM(27928) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(27928))))  severity failure;
	assert RAM(27929) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27929))))  severity failure;
	assert RAM(27930) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(27930))))  severity failure;
	assert RAM(27931) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(27931))))  severity failure;
	assert RAM(27932) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(27932))))  severity failure;
	assert RAM(27933) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(27933))))  severity failure;
	assert RAM(27934) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(27934))))  severity failure;
	assert RAM(27935) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(27935))))  severity failure;
	assert RAM(27936) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(27936))))  severity failure;
	assert RAM(27937) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(27937))))  severity failure;
	assert RAM(27938) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(27938))))  severity failure;
	assert RAM(27939) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(27939))))  severity failure;
	assert RAM(27940) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(27940))))  severity failure;
	assert RAM(27941) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(27941))))  severity failure;
	assert RAM(27942) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27942))))  severity failure;
	assert RAM(27943) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(27943))))  severity failure;
	assert RAM(27944) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(27944))))  severity failure;
	assert RAM(27945) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(27945))))  severity failure;
	assert RAM(27946) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(27946))))  severity failure;
	assert RAM(27947) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(27947))))  severity failure;
	assert RAM(27948) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27948))))  severity failure;
	assert RAM(27949) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27949))))  severity failure;
	assert RAM(27950) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(27950))))  severity failure;
	assert RAM(27951) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(27951))))  severity failure;
	assert RAM(27952) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(27952))))  severity failure;
	assert RAM(27953) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(27953))))  severity failure;
	assert RAM(27954) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(27954))))  severity failure;
	assert RAM(27955) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(27955))))  severity failure;
	assert RAM(27956) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(27956))))  severity failure;
	assert RAM(27957) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(27957))))  severity failure;
	assert RAM(27958) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(27958))))  severity failure;
	assert RAM(27959) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(27959))))  severity failure;
	assert RAM(27960) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(27960))))  severity failure;
	assert RAM(27961) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(27961))))  severity failure;
	assert RAM(27962) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(27962))))  severity failure;
	assert RAM(27963) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(27963))))  severity failure;
	assert RAM(27964) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(27964))))  severity failure;
	assert RAM(27965) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(27965))))  severity failure;
	assert RAM(27966) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(27966))))  severity failure;
	assert RAM(27967) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(27967))))  severity failure;
	assert RAM(27968) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(27968))))  severity failure;
	assert RAM(27969) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(27969))))  severity failure;
	assert RAM(27970) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(27970))))  severity failure;
	assert RAM(27971) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(27971))))  severity failure;
	assert RAM(27972) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(27972))))  severity failure;
	assert RAM(27973) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(27973))))  severity failure;
	assert RAM(27974) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(27974))))  severity failure;
	assert RAM(27975) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(27975))))  severity failure;
	assert RAM(27976) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(27976))))  severity failure;
	assert RAM(27977) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(27977))))  severity failure;
	assert RAM(27978) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(27978))))  severity failure;
	assert RAM(27979) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(27979))))  severity failure;
	assert RAM(27980) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(27980))))  severity failure;
	assert RAM(27981) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(27981))))  severity failure;
	assert RAM(27982) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(27982))))  severity failure;
	assert RAM(27983) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(27983))))  severity failure;
	assert RAM(27984) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(27984))))  severity failure;
	assert RAM(27985) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(27985))))  severity failure;
	assert RAM(27986) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(27986))))  severity failure;
	assert RAM(27987) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(27987))))  severity failure;
	assert RAM(27988) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(27988))))  severity failure;
	assert RAM(27989) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(27989))))  severity failure;
	assert RAM(27990) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(27990))))  severity failure;
	assert RAM(27991) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(27991))))  severity failure;
	assert RAM(27992) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(27992))))  severity failure;
	assert RAM(27993) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(27993))))  severity failure;
	assert RAM(27994) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(27994))))  severity failure;
	assert RAM(27995) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(27995))))  severity failure;
	assert RAM(27996) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(27996))))  severity failure;
	assert RAM(27997) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(27997))))  severity failure;
	assert RAM(27998) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(27998))))  severity failure;
	assert RAM(27999) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(27999))))  severity failure;
	assert RAM(28000) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28000))))  severity failure;
	assert RAM(28001) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(28001))))  severity failure;
	assert RAM(28002) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(28002))))  severity failure;
	assert RAM(28003) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(28003))))  severity failure;
	assert RAM(28004) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28004))))  severity failure;
	assert RAM(28005) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(28005))))  severity failure;
	assert RAM(28006) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(28006))))  severity failure;
	assert RAM(28007) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28007))))  severity failure;
	assert RAM(28008) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(28008))))  severity failure;
	assert RAM(28009) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(28009))))  severity failure;
	assert RAM(28010) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(28010))))  severity failure;
	assert RAM(28011) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28011))))  severity failure;
	assert RAM(28012) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(28012))))  severity failure;
	assert RAM(28013) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28013))))  severity failure;
	assert RAM(28014) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(28014))))  severity failure;
	assert RAM(28015) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28015))))  severity failure;
	assert RAM(28016) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(28016))))  severity failure;
	assert RAM(28017) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28017))))  severity failure;
	assert RAM(28018) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(28018))))  severity failure;
	assert RAM(28019) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(28019))))  severity failure;
	assert RAM(28020) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(28020))))  severity failure;
	assert RAM(28021) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(28021))))  severity failure;
	assert RAM(28022) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28022))))  severity failure;
	assert RAM(28023) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(28023))))  severity failure;
	assert RAM(28024) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28024))))  severity failure;
	assert RAM(28025) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(28025))))  severity failure;
	assert RAM(28026) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28026))))  severity failure;
	assert RAM(28027) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(28027))))  severity failure;
	assert RAM(28028) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28028))))  severity failure;
	assert RAM(28029) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28029))))  severity failure;
	assert RAM(28030) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(28030))))  severity failure;
	assert RAM(28031) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28031))))  severity failure;
	assert RAM(28032) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(28032))))  severity failure;
	assert RAM(28033) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(28033))))  severity failure;
	assert RAM(28034) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(28034))))  severity failure;
	assert RAM(28035) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28035))))  severity failure;
	assert RAM(28036) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28036))))  severity failure;
	assert RAM(28037) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28037))))  severity failure;
	assert RAM(28038) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28038))))  severity failure;
	assert RAM(28039) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28039))))  severity failure;
	assert RAM(28040) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(28040))))  severity failure;
	assert RAM(28041) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28041))))  severity failure;
	assert RAM(28042) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28042))))  severity failure;
	assert RAM(28043) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28043))))  severity failure;
	assert RAM(28044) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(28044))))  severity failure;
	assert RAM(28045) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(28045))))  severity failure;
	assert RAM(28046) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28046))))  severity failure;
	assert RAM(28047) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(28047))))  severity failure;
	assert RAM(28048) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(28048))))  severity failure;
	assert RAM(28049) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(28049))))  severity failure;
	assert RAM(28050) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28050))))  severity failure;
	assert RAM(28051) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(28051))))  severity failure;
	assert RAM(28052) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(28052))))  severity failure;
	assert RAM(28053) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(28053))))  severity failure;
	assert RAM(28054) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28054))))  severity failure;
	assert RAM(28055) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28055))))  severity failure;
	assert RAM(28056) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(28056))))  severity failure;
	assert RAM(28057) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(28057))))  severity failure;
	assert RAM(28058) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(28058))))  severity failure;
	assert RAM(28059) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(28059))))  severity failure;
	assert RAM(28060) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28060))))  severity failure;
	assert RAM(28061) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(28061))))  severity failure;
	assert RAM(28062) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28062))))  severity failure;
	assert RAM(28063) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28063))))  severity failure;
	assert RAM(28064) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(28064))))  severity failure;
	assert RAM(28065) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(28065))))  severity failure;
	assert RAM(28066) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(28066))))  severity failure;
	assert RAM(28067) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(28067))))  severity failure;
	assert RAM(28068) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28068))))  severity failure;
	assert RAM(28069) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(28069))))  severity failure;
	assert RAM(28070) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(28070))))  severity failure;
	assert RAM(28071) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28071))))  severity failure;
	assert RAM(28072) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(28072))))  severity failure;
	assert RAM(28073) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28073))))  severity failure;
	assert RAM(28074) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(28074))))  severity failure;
	assert RAM(28075) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28075))))  severity failure;
	assert RAM(28076) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28076))))  severity failure;
	assert RAM(28077) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(28077))))  severity failure;
	assert RAM(28078) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(28078))))  severity failure;
	assert RAM(28079) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(28079))))  severity failure;
	assert RAM(28080) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(28080))))  severity failure;
	assert RAM(28081) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28081))))  severity failure;
	assert RAM(28082) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(28082))))  severity failure;
	assert RAM(28083) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(28083))))  severity failure;
	assert RAM(28084) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(28084))))  severity failure;
	assert RAM(28085) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(28085))))  severity failure;
	assert RAM(28086) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28086))))  severity failure;
	assert RAM(28087) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(28087))))  severity failure;
	assert RAM(28088) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28088))))  severity failure;
	assert RAM(28089) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(28089))))  severity failure;
	assert RAM(28090) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(28090))))  severity failure;
	assert RAM(28091) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(28091))))  severity failure;
	assert RAM(28092) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(28092))))  severity failure;
	assert RAM(28093) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28093))))  severity failure;
	assert RAM(28094) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(28094))))  severity failure;
	assert RAM(28095) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(28095))))  severity failure;
	assert RAM(28096) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(28096))))  severity failure;
	assert RAM(28097) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28097))))  severity failure;
	assert RAM(28098) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28098))))  severity failure;
	assert RAM(28099) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28099))))  severity failure;
	assert RAM(28100) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28100))))  severity failure;
	assert RAM(28101) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(28101))))  severity failure;
	assert RAM(28102) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(28102))))  severity failure;
	assert RAM(28103) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28103))))  severity failure;
	assert RAM(28104) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28104))))  severity failure;
	assert RAM(28105) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(28105))))  severity failure;
	assert RAM(28106) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(28106))))  severity failure;
	assert RAM(28107) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(28107))))  severity failure;
	assert RAM(28108) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(28108))))  severity failure;
	assert RAM(28109) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(28109))))  severity failure;
	assert RAM(28110) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28110))))  severity failure;
	assert RAM(28111) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(28111))))  severity failure;
	assert RAM(28112) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(28112))))  severity failure;
	assert RAM(28113) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(28113))))  severity failure;
	assert RAM(28114) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28114))))  severity failure;
	assert RAM(28115) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(28115))))  severity failure;
	assert RAM(28116) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(28116))))  severity failure;
	assert RAM(28117) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(28117))))  severity failure;
	assert RAM(28118) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(28118))))  severity failure;
	assert RAM(28119) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28119))))  severity failure;
	assert RAM(28120) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(28120))))  severity failure;
	assert RAM(28121) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28121))))  severity failure;
	assert RAM(28122) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(28122))))  severity failure;
	assert RAM(28123) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(28123))))  severity failure;
	assert RAM(28124) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28124))))  severity failure;
	assert RAM(28125) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28125))))  severity failure;
	assert RAM(28126) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(28126))))  severity failure;
	assert RAM(28127) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(28127))))  severity failure;
	assert RAM(28128) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(28128))))  severity failure;
	assert RAM(28129) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(28129))))  severity failure;
	assert RAM(28130) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(28130))))  severity failure;
	assert RAM(28131) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(28131))))  severity failure;
	assert RAM(28132) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(28132))))  severity failure;
	assert RAM(28133) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(28133))))  severity failure;
	assert RAM(28134) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28134))))  severity failure;
	assert RAM(28135) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(28135))))  severity failure;
	assert RAM(28136) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28136))))  severity failure;
	assert RAM(28137) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(28137))))  severity failure;
	assert RAM(28138) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(28138))))  severity failure;
	assert RAM(28139) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28139))))  severity failure;
	assert RAM(28140) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(28140))))  severity failure;
	assert RAM(28141) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28141))))  severity failure;
	assert RAM(28142) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(28142))))  severity failure;
	assert RAM(28143) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(28143))))  severity failure;
	assert RAM(28144) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28144))))  severity failure;
	assert RAM(28145) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(28145))))  severity failure;
	assert RAM(28146) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28146))))  severity failure;
	assert RAM(28147) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28147))))  severity failure;
	assert RAM(28148) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(28148))))  severity failure;
	assert RAM(28149) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(28149))))  severity failure;
	assert RAM(28150) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28150))))  severity failure;
	assert RAM(28151) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28151))))  severity failure;
	assert RAM(28152) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(28152))))  severity failure;
	assert RAM(28153) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(28153))))  severity failure;
	assert RAM(28154) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(28154))))  severity failure;
	assert RAM(28155) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28155))))  severity failure;
	assert RAM(28156) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(28156))))  severity failure;
	assert RAM(28157) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28157))))  severity failure;
	assert RAM(28158) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28158))))  severity failure;
	assert RAM(28159) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28159))))  severity failure;
	assert RAM(28160) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28160))))  severity failure;
	assert RAM(28161) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28161))))  severity failure;
	assert RAM(28162) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28162))))  severity failure;
	assert RAM(28163) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(28163))))  severity failure;
	assert RAM(28164) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(28164))))  severity failure;
	assert RAM(28165) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(28165))))  severity failure;
	assert RAM(28166) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28166))))  severity failure;
	assert RAM(28167) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(28167))))  severity failure;
	assert RAM(28168) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(28168))))  severity failure;
	assert RAM(28169) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28169))))  severity failure;
	assert RAM(28170) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(28170))))  severity failure;
	assert RAM(28171) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(28171))))  severity failure;
	assert RAM(28172) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(28172))))  severity failure;
	assert RAM(28173) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(28173))))  severity failure;
	assert RAM(28174) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(28174))))  severity failure;
	assert RAM(28175) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28175))))  severity failure;
	assert RAM(28176) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28176))))  severity failure;
	assert RAM(28177) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(28177))))  severity failure;
	assert RAM(28178) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(28178))))  severity failure;
	assert RAM(28179) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(28179))))  severity failure;
	assert RAM(28180) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(28180))))  severity failure;
	assert RAM(28181) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(28181))))  severity failure;
	assert RAM(28182) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(28182))))  severity failure;
	assert RAM(28183) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(28183))))  severity failure;
	assert RAM(28184) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28184))))  severity failure;
	assert RAM(28185) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28185))))  severity failure;
	assert RAM(28186) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28186))))  severity failure;
	assert RAM(28187) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28187))))  severity failure;
	assert RAM(28188) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(28188))))  severity failure;
	assert RAM(28189) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28189))))  severity failure;
	assert RAM(28190) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28190))))  severity failure;
	assert RAM(28191) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(28191))))  severity failure;
	assert RAM(28192) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(28192))))  severity failure;
	assert RAM(28193) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(28193))))  severity failure;
	assert RAM(28194) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28194))))  severity failure;
	assert RAM(28195) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(28195))))  severity failure;
	assert RAM(28196) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(28196))))  severity failure;
	assert RAM(28197) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(28197))))  severity failure;
	assert RAM(28198) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28198))))  severity failure;
	assert RAM(28199) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(28199))))  severity failure;
	assert RAM(28200) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(28200))))  severity failure;
	assert RAM(28201) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(28201))))  severity failure;
	assert RAM(28202) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28202))))  severity failure;
	assert RAM(28203) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(28203))))  severity failure;
	assert RAM(28204) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28204))))  severity failure;
	assert RAM(28205) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(28205))))  severity failure;
	assert RAM(28206) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(28206))))  severity failure;
	assert RAM(28207) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28207))))  severity failure;
	assert RAM(28208) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(28208))))  severity failure;
	assert RAM(28209) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28209))))  severity failure;
	assert RAM(28210) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(28210))))  severity failure;
	assert RAM(28211) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(28211))))  severity failure;
	assert RAM(28212) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(28212))))  severity failure;
	assert RAM(28213) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(28213))))  severity failure;
	assert RAM(28214) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(28214))))  severity failure;
	assert RAM(28215) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(28215))))  severity failure;
	assert RAM(28216) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(28216))))  severity failure;
	assert RAM(28217) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28217))))  severity failure;
	assert RAM(28218) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(28218))))  severity failure;
	assert RAM(28219) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28219))))  severity failure;
	assert RAM(28220) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28220))))  severity failure;
	assert RAM(28221) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28221))))  severity failure;
	assert RAM(28222) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(28222))))  severity failure;
	assert RAM(28223) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28223))))  severity failure;
	assert RAM(28224) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(28224))))  severity failure;
	assert RAM(28225) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(28225))))  severity failure;
	assert RAM(28226) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(28226))))  severity failure;
	assert RAM(28227) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28227))))  severity failure;
	assert RAM(28228) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(28228))))  severity failure;
	assert RAM(28229) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(28229))))  severity failure;
	assert RAM(28230) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(28230))))  severity failure;
	assert RAM(28231) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(28231))))  severity failure;
	assert RAM(28232) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(28232))))  severity failure;
	assert RAM(28233) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(28233))))  severity failure;
	assert RAM(28234) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(28234))))  severity failure;
	assert RAM(28235) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(28235))))  severity failure;
	assert RAM(28236) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(28236))))  severity failure;
	assert RAM(28237) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(28237))))  severity failure;
	assert RAM(28238) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(28238))))  severity failure;
	assert RAM(28239) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(28239))))  severity failure;
	assert RAM(28240) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28240))))  severity failure;
	assert RAM(28241) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(28241))))  severity failure;
	assert RAM(28242) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(28242))))  severity failure;
	assert RAM(28243) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(28243))))  severity failure;
	assert RAM(28244) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28244))))  severity failure;
	assert RAM(28245) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28245))))  severity failure;
	assert RAM(28246) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(28246))))  severity failure;
	assert RAM(28247) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28247))))  severity failure;
	assert RAM(28248) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(28248))))  severity failure;
	assert RAM(28249) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(28249))))  severity failure;
	assert RAM(28250) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(28250))))  severity failure;
	assert RAM(28251) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28251))))  severity failure;
	assert RAM(28252) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(28252))))  severity failure;
	assert RAM(28253) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(28253))))  severity failure;
	assert RAM(28254) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(28254))))  severity failure;
	assert RAM(28255) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28255))))  severity failure;
	assert RAM(28256) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(28256))))  severity failure;
	assert RAM(28257) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28257))))  severity failure;
	assert RAM(28258) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(28258))))  severity failure;
	assert RAM(28259) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(28259))))  severity failure;
	assert RAM(28260) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28260))))  severity failure;
	assert RAM(28261) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28261))))  severity failure;
	assert RAM(28262) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(28262))))  severity failure;
	assert RAM(28263) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28263))))  severity failure;
	assert RAM(28264) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(28264))))  severity failure;
	assert RAM(28265) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(28265))))  severity failure;
	assert RAM(28266) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28266))))  severity failure;
	assert RAM(28267) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(28267))))  severity failure;
	assert RAM(28268) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(28268))))  severity failure;
	assert RAM(28269) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(28269))))  severity failure;
	assert RAM(28270) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(28270))))  severity failure;
	assert RAM(28271) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(28271))))  severity failure;
	assert RAM(28272) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(28272))))  severity failure;
	assert RAM(28273) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28273))))  severity failure;
	assert RAM(28274) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(28274))))  severity failure;
	assert RAM(28275) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(28275))))  severity failure;
	assert RAM(28276) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(28276))))  severity failure;
	assert RAM(28277) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(28277))))  severity failure;
	assert RAM(28278) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28278))))  severity failure;
	assert RAM(28279) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28279))))  severity failure;
	assert RAM(28280) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(28280))))  severity failure;
	assert RAM(28281) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28281))))  severity failure;
	assert RAM(28282) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(28282))))  severity failure;
	assert RAM(28283) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(28283))))  severity failure;
	assert RAM(28284) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(28284))))  severity failure;
	assert RAM(28285) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(28285))))  severity failure;
	assert RAM(28286) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(28286))))  severity failure;
	assert RAM(28287) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(28287))))  severity failure;
	assert RAM(28288) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(28288))))  severity failure;
	assert RAM(28289) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28289))))  severity failure;
	assert RAM(28290) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28290))))  severity failure;
	assert RAM(28291) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(28291))))  severity failure;
	assert RAM(28292) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28292))))  severity failure;
	assert RAM(28293) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(28293))))  severity failure;
	assert RAM(28294) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(28294))))  severity failure;
	assert RAM(28295) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28295))))  severity failure;
	assert RAM(28296) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(28296))))  severity failure;
	assert RAM(28297) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28297))))  severity failure;
	assert RAM(28298) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28298))))  severity failure;
	assert RAM(28299) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(28299))))  severity failure;
	assert RAM(28300) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(28300))))  severity failure;
	assert RAM(28301) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(28301))))  severity failure;
	assert RAM(28302) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(28302))))  severity failure;
	assert RAM(28303) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28303))))  severity failure;
	assert RAM(28304) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(28304))))  severity failure;
	assert RAM(28305) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28305))))  severity failure;
	assert RAM(28306) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(28306))))  severity failure;
	assert RAM(28307) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28307))))  severity failure;
	assert RAM(28308) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(28308))))  severity failure;
	assert RAM(28309) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(28309))))  severity failure;
	assert RAM(28310) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(28310))))  severity failure;
	assert RAM(28311) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28311))))  severity failure;
	assert RAM(28312) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28312))))  severity failure;
	assert RAM(28313) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28313))))  severity failure;
	assert RAM(28314) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(28314))))  severity failure;
	assert RAM(28315) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(28315))))  severity failure;
	assert RAM(28316) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(28316))))  severity failure;
	assert RAM(28317) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(28317))))  severity failure;
	assert RAM(28318) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28318))))  severity failure;
	assert RAM(28319) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(28319))))  severity failure;
	assert RAM(28320) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28320))))  severity failure;
	assert RAM(28321) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(28321))))  severity failure;
	assert RAM(28322) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(28322))))  severity failure;
	assert RAM(28323) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(28323))))  severity failure;
	assert RAM(28324) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28324))))  severity failure;
	assert RAM(28325) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(28325))))  severity failure;
	assert RAM(28326) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(28326))))  severity failure;
	assert RAM(28327) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(28327))))  severity failure;
	assert RAM(28328) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28328))))  severity failure;
	assert RAM(28329) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(28329))))  severity failure;
	assert RAM(28330) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28330))))  severity failure;
	assert RAM(28331) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(28331))))  severity failure;
	assert RAM(28332) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(28332))))  severity failure;
	assert RAM(28333) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(28333))))  severity failure;
	assert RAM(28334) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28334))))  severity failure;
	assert RAM(28335) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(28335))))  severity failure;
	assert RAM(28336) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28336))))  severity failure;
	assert RAM(28337) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(28337))))  severity failure;
	assert RAM(28338) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28338))))  severity failure;
	assert RAM(28339) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(28339))))  severity failure;
	assert RAM(28340) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(28340))))  severity failure;
	assert RAM(28341) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(28341))))  severity failure;
	assert RAM(28342) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(28342))))  severity failure;
	assert RAM(28343) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(28343))))  severity failure;
	assert RAM(28344) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(28344))))  severity failure;
	assert RAM(28345) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28345))))  severity failure;
	assert RAM(28346) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(28346))))  severity failure;
	assert RAM(28347) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28347))))  severity failure;
	assert RAM(28348) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(28348))))  severity failure;
	assert RAM(28349) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28349))))  severity failure;
	assert RAM(28350) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(28350))))  severity failure;
	assert RAM(28351) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(28351))))  severity failure;
	assert RAM(28352) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(28352))))  severity failure;
	assert RAM(28353) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28353))))  severity failure;
	assert RAM(28354) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28354))))  severity failure;
	assert RAM(28355) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28355))))  severity failure;
	assert RAM(28356) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28356))))  severity failure;
	assert RAM(28357) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(28357))))  severity failure;
	assert RAM(28358) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28358))))  severity failure;
	assert RAM(28359) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(28359))))  severity failure;
	assert RAM(28360) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(28360))))  severity failure;
	assert RAM(28361) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28361))))  severity failure;
	assert RAM(28362) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(28362))))  severity failure;
	assert RAM(28363) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(28363))))  severity failure;
	assert RAM(28364) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(28364))))  severity failure;
	assert RAM(28365) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(28365))))  severity failure;
	assert RAM(28366) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(28366))))  severity failure;
	assert RAM(28367) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(28367))))  severity failure;
	assert RAM(28368) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(28368))))  severity failure;
	assert RAM(28369) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28369))))  severity failure;
	assert RAM(28370) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(28370))))  severity failure;
	assert RAM(28371) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(28371))))  severity failure;
	assert RAM(28372) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28372))))  severity failure;
	assert RAM(28373) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(28373))))  severity failure;
	assert RAM(28374) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(28374))))  severity failure;
	assert RAM(28375) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28375))))  severity failure;
	assert RAM(28376) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28376))))  severity failure;
	assert RAM(28377) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28377))))  severity failure;
	assert RAM(28378) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(28378))))  severity failure;
	assert RAM(28379) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(28379))))  severity failure;
	assert RAM(28380) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(28380))))  severity failure;
	assert RAM(28381) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28381))))  severity failure;
	assert RAM(28382) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28382))))  severity failure;
	assert RAM(28383) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(28383))))  severity failure;
	assert RAM(28384) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(28384))))  severity failure;
	assert RAM(28385) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(28385))))  severity failure;
	assert RAM(28386) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28386))))  severity failure;
	assert RAM(28387) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28387))))  severity failure;
	assert RAM(28388) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28388))))  severity failure;
	assert RAM(28389) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28389))))  severity failure;
	assert RAM(28390) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28390))))  severity failure;
	assert RAM(28391) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(28391))))  severity failure;
	assert RAM(28392) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(28392))))  severity failure;
	assert RAM(28393) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(28393))))  severity failure;
	assert RAM(28394) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28394))))  severity failure;
	assert RAM(28395) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28395))))  severity failure;
	assert RAM(28396) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28396))))  severity failure;
	assert RAM(28397) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(28397))))  severity failure;
	assert RAM(28398) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28398))))  severity failure;
	assert RAM(28399) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(28399))))  severity failure;
	assert RAM(28400) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(28400))))  severity failure;
	assert RAM(28401) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(28401))))  severity failure;
	assert RAM(28402) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(28402))))  severity failure;
	assert RAM(28403) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(28403))))  severity failure;
	assert RAM(28404) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(28404))))  severity failure;
	assert RAM(28405) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(28405))))  severity failure;
	assert RAM(28406) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(28406))))  severity failure;
	assert RAM(28407) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(28407))))  severity failure;
	assert RAM(28408) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(28408))))  severity failure;
	assert RAM(28409) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(28409))))  severity failure;
	assert RAM(28410) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(28410))))  severity failure;
	assert RAM(28411) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(28411))))  severity failure;
	assert RAM(28412) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(28412))))  severity failure;
	assert RAM(28413) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(28413))))  severity failure;
	assert RAM(28414) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(28414))))  severity failure;
	assert RAM(28415) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(28415))))  severity failure;
	assert RAM(28416) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(28416))))  severity failure;
	assert RAM(28417) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(28417))))  severity failure;
	assert RAM(28418) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(28418))))  severity failure;
	assert RAM(28419) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28419))))  severity failure;
	assert RAM(28420) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(28420))))  severity failure;
	assert RAM(28421) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(28421))))  severity failure;
	assert RAM(28422) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(28422))))  severity failure;
	assert RAM(28423) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(28423))))  severity failure;
	assert RAM(28424) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(28424))))  severity failure;
	assert RAM(28425) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(28425))))  severity failure;
	assert RAM(28426) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(28426))))  severity failure;
	assert RAM(28427) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(28427))))  severity failure;
	assert RAM(28428) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28428))))  severity failure;
	assert RAM(28429) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28429))))  severity failure;
	assert RAM(28430) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(28430))))  severity failure;
	assert RAM(28431) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28431))))  severity failure;
	assert RAM(28432) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(28432))))  severity failure;
	assert RAM(28433) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(28433))))  severity failure;
	assert RAM(28434) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(28434))))  severity failure;
	assert RAM(28435) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28435))))  severity failure;
	assert RAM(28436) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(28436))))  severity failure;
	assert RAM(28437) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28437))))  severity failure;
	assert RAM(28438) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(28438))))  severity failure;
	assert RAM(28439) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(28439))))  severity failure;
	assert RAM(28440) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28440))))  severity failure;
	assert RAM(28441) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(28441))))  severity failure;
	assert RAM(28442) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(28442))))  severity failure;
	assert RAM(28443) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28443))))  severity failure;
	assert RAM(28444) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(28444))))  severity failure;
	assert RAM(28445) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(28445))))  severity failure;
	assert RAM(28446) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28446))))  severity failure;
	assert RAM(28447) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28447))))  severity failure;
	assert RAM(28448) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(28448))))  severity failure;
	assert RAM(28449) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(28449))))  severity failure;
	assert RAM(28450) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28450))))  severity failure;
	assert RAM(28451) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28451))))  severity failure;
	assert RAM(28452) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(28452))))  severity failure;
	assert RAM(28453) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28453))))  severity failure;
	assert RAM(28454) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(28454))))  severity failure;
	assert RAM(28455) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(28455))))  severity failure;
	assert RAM(28456) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(28456))))  severity failure;
	assert RAM(28457) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28457))))  severity failure;
	assert RAM(28458) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(28458))))  severity failure;
	assert RAM(28459) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(28459))))  severity failure;
	assert RAM(28460) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(28460))))  severity failure;
	assert RAM(28461) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28461))))  severity failure;
	assert RAM(28462) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(28462))))  severity failure;
	assert RAM(28463) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28463))))  severity failure;
	assert RAM(28464) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(28464))))  severity failure;
	assert RAM(28465) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(28465))))  severity failure;
	assert RAM(28466) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(28466))))  severity failure;
	assert RAM(28467) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(28467))))  severity failure;
	assert RAM(28468) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(28468))))  severity failure;
	assert RAM(28469) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(28469))))  severity failure;
	assert RAM(28470) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(28470))))  severity failure;
	assert RAM(28471) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(28471))))  severity failure;
	assert RAM(28472) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(28472))))  severity failure;
	assert RAM(28473) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(28473))))  severity failure;
	assert RAM(28474) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(28474))))  severity failure;
	assert RAM(28475) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28475))))  severity failure;
	assert RAM(28476) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(28476))))  severity failure;
	assert RAM(28477) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(28477))))  severity failure;
	assert RAM(28478) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(28478))))  severity failure;
	assert RAM(28479) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(28479))))  severity failure;
	assert RAM(28480) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(28480))))  severity failure;
	assert RAM(28481) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(28481))))  severity failure;
	assert RAM(28482) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28482))))  severity failure;
	assert RAM(28483) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28483))))  severity failure;
	assert RAM(28484) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(28484))))  severity failure;
	assert RAM(28485) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(28485))))  severity failure;
	assert RAM(28486) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(28486))))  severity failure;
	assert RAM(28487) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(28487))))  severity failure;
	assert RAM(28488) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(28488))))  severity failure;
	assert RAM(28489) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28489))))  severity failure;
	assert RAM(28490) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(28490))))  severity failure;
	assert RAM(28491) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(28491))))  severity failure;
	assert RAM(28492) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(28492))))  severity failure;
	assert RAM(28493) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(28493))))  severity failure;
	assert RAM(28494) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(28494))))  severity failure;
	assert RAM(28495) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28495))))  severity failure;
	assert RAM(28496) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(28496))))  severity failure;
	assert RAM(28497) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(28497))))  severity failure;
	assert RAM(28498) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(28498))))  severity failure;
	assert RAM(28499) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28499))))  severity failure;
	assert RAM(28500) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28500))))  severity failure;
	assert RAM(28501) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(28501))))  severity failure;
	assert RAM(28502) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28502))))  severity failure;
	assert RAM(28503) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(28503))))  severity failure;
	assert RAM(28504) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(28504))))  severity failure;
	assert RAM(28505) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(28505))))  severity failure;
	assert RAM(28506) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(28506))))  severity failure;
	assert RAM(28507) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28507))))  severity failure;
	assert RAM(28508) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28508))))  severity failure;
	assert RAM(28509) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(28509))))  severity failure;
	assert RAM(28510) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(28510))))  severity failure;
	assert RAM(28511) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(28511))))  severity failure;
	assert RAM(28512) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28512))))  severity failure;
	assert RAM(28513) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(28513))))  severity failure;
	assert RAM(28514) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(28514))))  severity failure;
	assert RAM(28515) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28515))))  severity failure;
	assert RAM(28516) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28516))))  severity failure;
	assert RAM(28517) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28517))))  severity failure;
	assert RAM(28518) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28518))))  severity failure;
	assert RAM(28519) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(28519))))  severity failure;
	assert RAM(28520) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(28520))))  severity failure;
	assert RAM(28521) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(28521))))  severity failure;
	assert RAM(28522) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28522))))  severity failure;
	assert RAM(28523) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(28523))))  severity failure;
	assert RAM(28524) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(28524))))  severity failure;
	assert RAM(28525) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28525))))  severity failure;
	assert RAM(28526) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28526))))  severity failure;
	assert RAM(28527) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(28527))))  severity failure;
	assert RAM(28528) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28528))))  severity failure;
	assert RAM(28529) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28529))))  severity failure;
	assert RAM(28530) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(28530))))  severity failure;
	assert RAM(28531) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(28531))))  severity failure;
	assert RAM(28532) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(28532))))  severity failure;
	assert RAM(28533) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28533))))  severity failure;
	assert RAM(28534) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(28534))))  severity failure;
	assert RAM(28535) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(28535))))  severity failure;
	assert RAM(28536) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28536))))  severity failure;
	assert RAM(28537) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(28537))))  severity failure;
	assert RAM(28538) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(28538))))  severity failure;
	assert RAM(28539) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28539))))  severity failure;
	assert RAM(28540) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(28540))))  severity failure;
	assert RAM(28541) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28541))))  severity failure;
	assert RAM(28542) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(28542))))  severity failure;
	assert RAM(28543) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(28543))))  severity failure;
	assert RAM(28544) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(28544))))  severity failure;
	assert RAM(28545) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(28545))))  severity failure;
	assert RAM(28546) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(28546))))  severity failure;
	assert RAM(28547) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28547))))  severity failure;
	assert RAM(28548) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(28548))))  severity failure;
	assert RAM(28549) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28549))))  severity failure;
	assert RAM(28550) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(28550))))  severity failure;
	assert RAM(28551) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28551))))  severity failure;
	assert RAM(28552) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(28552))))  severity failure;
	assert RAM(28553) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28553))))  severity failure;
	assert RAM(28554) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(28554))))  severity failure;
	assert RAM(28555) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(28555))))  severity failure;
	assert RAM(28556) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(28556))))  severity failure;
	assert RAM(28557) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(28557))))  severity failure;
	assert RAM(28558) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28558))))  severity failure;
	assert RAM(28559) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(28559))))  severity failure;
	assert RAM(28560) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28560))))  severity failure;
	assert RAM(28561) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(28561))))  severity failure;
	assert RAM(28562) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(28562))))  severity failure;
	assert RAM(28563) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28563))))  severity failure;
	assert RAM(28564) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(28564))))  severity failure;
	assert RAM(28565) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(28565))))  severity failure;
	assert RAM(28566) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28566))))  severity failure;
	assert RAM(28567) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(28567))))  severity failure;
	assert RAM(28568) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(28568))))  severity failure;
	assert RAM(28569) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(28569))))  severity failure;
	assert RAM(28570) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(28570))))  severity failure;
	assert RAM(28571) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28571))))  severity failure;
	assert RAM(28572) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(28572))))  severity failure;
	assert RAM(28573) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(28573))))  severity failure;
	assert RAM(28574) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(28574))))  severity failure;
	assert RAM(28575) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(28575))))  severity failure;
	assert RAM(28576) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28576))))  severity failure;
	assert RAM(28577) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28577))))  severity failure;
	assert RAM(28578) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(28578))))  severity failure;
	assert RAM(28579) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28579))))  severity failure;
	assert RAM(28580) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28580))))  severity failure;
	assert RAM(28581) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(28581))))  severity failure;
	assert RAM(28582) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(28582))))  severity failure;
	assert RAM(28583) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(28583))))  severity failure;
	assert RAM(28584) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(28584))))  severity failure;
	assert RAM(28585) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(28585))))  severity failure;
	assert RAM(28586) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28586))))  severity failure;
	assert RAM(28587) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(28587))))  severity failure;
	assert RAM(28588) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(28588))))  severity failure;
	assert RAM(28589) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28589))))  severity failure;
	assert RAM(28590) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28590))))  severity failure;
	assert RAM(28591) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28591))))  severity failure;
	assert RAM(28592) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(28592))))  severity failure;
	assert RAM(28593) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28593))))  severity failure;
	assert RAM(28594) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(28594))))  severity failure;
	assert RAM(28595) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(28595))))  severity failure;
	assert RAM(28596) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28596))))  severity failure;
	assert RAM(28597) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28597))))  severity failure;
	assert RAM(28598) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(28598))))  severity failure;
	assert RAM(28599) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28599))))  severity failure;
	assert RAM(28600) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(28600))))  severity failure;
	assert RAM(28601) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(28601))))  severity failure;
	assert RAM(28602) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(28602))))  severity failure;
	assert RAM(28603) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(28603))))  severity failure;
	assert RAM(28604) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(28604))))  severity failure;
	assert RAM(28605) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(28605))))  severity failure;
	assert RAM(28606) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(28606))))  severity failure;
	assert RAM(28607) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(28607))))  severity failure;
	assert RAM(28608) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(28608))))  severity failure;
	assert RAM(28609) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(28609))))  severity failure;
	assert RAM(28610) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(28610))))  severity failure;
	assert RAM(28611) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(28611))))  severity failure;
	assert RAM(28612) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28612))))  severity failure;
	assert RAM(28613) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28613))))  severity failure;
	assert RAM(28614) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(28614))))  severity failure;
	assert RAM(28615) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(28615))))  severity failure;
	assert RAM(28616) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28616))))  severity failure;
	assert RAM(28617) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(28617))))  severity failure;
	assert RAM(28618) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(28618))))  severity failure;
	assert RAM(28619) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28619))))  severity failure;
	assert RAM(28620) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(28620))))  severity failure;
	assert RAM(28621) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(28621))))  severity failure;
	assert RAM(28622) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(28622))))  severity failure;
	assert RAM(28623) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28623))))  severity failure;
	assert RAM(28624) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(28624))))  severity failure;
	assert RAM(28625) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(28625))))  severity failure;
	assert RAM(28626) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(28626))))  severity failure;
	assert RAM(28627) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(28627))))  severity failure;
	assert RAM(28628) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(28628))))  severity failure;
	assert RAM(28629) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(28629))))  severity failure;
	assert RAM(28630) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(28630))))  severity failure;
	assert RAM(28631) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(28631))))  severity failure;
	assert RAM(28632) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28632))))  severity failure;
	assert RAM(28633) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28633))))  severity failure;
	assert RAM(28634) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28634))))  severity failure;
	assert RAM(28635) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28635))))  severity failure;
	assert RAM(28636) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(28636))))  severity failure;
	assert RAM(28637) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(28637))))  severity failure;
	assert RAM(28638) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(28638))))  severity failure;
	assert RAM(28639) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28639))))  severity failure;
	assert RAM(28640) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(28640))))  severity failure;
	assert RAM(28641) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(28641))))  severity failure;
	assert RAM(28642) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(28642))))  severity failure;
	assert RAM(28643) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(28643))))  severity failure;
	assert RAM(28644) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(28644))))  severity failure;
	assert RAM(28645) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28645))))  severity failure;
	assert RAM(28646) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28646))))  severity failure;
	assert RAM(28647) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(28647))))  severity failure;
	assert RAM(28648) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(28648))))  severity failure;
	assert RAM(28649) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(28649))))  severity failure;
	assert RAM(28650) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28650))))  severity failure;
	assert RAM(28651) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(28651))))  severity failure;
	assert RAM(28652) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28652))))  severity failure;
	assert RAM(28653) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(28653))))  severity failure;
	assert RAM(28654) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(28654))))  severity failure;
	assert RAM(28655) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(28655))))  severity failure;
	assert RAM(28656) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(28656))))  severity failure;
	assert RAM(28657) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(28657))))  severity failure;
	assert RAM(28658) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28658))))  severity failure;
	assert RAM(28659) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(28659))))  severity failure;
	assert RAM(28660) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28660))))  severity failure;
	assert RAM(28661) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(28661))))  severity failure;
	assert RAM(28662) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(28662))))  severity failure;
	assert RAM(28663) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28663))))  severity failure;
	assert RAM(28664) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28664))))  severity failure;
	assert RAM(28665) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28665))))  severity failure;
	assert RAM(28666) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28666))))  severity failure;
	assert RAM(28667) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28667))))  severity failure;
	assert RAM(28668) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(28668))))  severity failure;
	assert RAM(28669) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(28669))))  severity failure;
	assert RAM(28670) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(28670))))  severity failure;
	assert RAM(28671) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(28671))))  severity failure;
	assert RAM(28672) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(28672))))  severity failure;
	assert RAM(28673) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(28673))))  severity failure;
	assert RAM(28674) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(28674))))  severity failure;
	assert RAM(28675) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28675))))  severity failure;
	assert RAM(28676) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(28676))))  severity failure;
	assert RAM(28677) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(28677))))  severity failure;
	assert RAM(28678) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(28678))))  severity failure;
	assert RAM(28679) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28679))))  severity failure;
	assert RAM(28680) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(28680))))  severity failure;
	assert RAM(28681) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(28681))))  severity failure;
	assert RAM(28682) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28682))))  severity failure;
	assert RAM(28683) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(28683))))  severity failure;
	assert RAM(28684) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(28684))))  severity failure;
	assert RAM(28685) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(28685))))  severity failure;
	assert RAM(28686) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(28686))))  severity failure;
	assert RAM(28687) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(28687))))  severity failure;
	assert RAM(28688) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(28688))))  severity failure;
	assert RAM(28689) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(28689))))  severity failure;
	assert RAM(28690) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(28690))))  severity failure;
	assert RAM(28691) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(28691))))  severity failure;
	assert RAM(28692) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(28692))))  severity failure;
	assert RAM(28693) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28693))))  severity failure;
	assert RAM(28694) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(28694))))  severity failure;
	assert RAM(28695) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(28695))))  severity failure;
	assert RAM(28696) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28696))))  severity failure;
	assert RAM(28697) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28697))))  severity failure;
	assert RAM(28698) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(28698))))  severity failure;
	assert RAM(28699) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28699))))  severity failure;
	assert RAM(28700) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(28700))))  severity failure;
	assert RAM(28701) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28701))))  severity failure;
	assert RAM(28702) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(28702))))  severity failure;
	assert RAM(28703) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(28703))))  severity failure;
	assert RAM(28704) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(28704))))  severity failure;
	assert RAM(28705) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(28705))))  severity failure;
	assert RAM(28706) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(28706))))  severity failure;
	assert RAM(28707) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(28707))))  severity failure;
	assert RAM(28708) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28708))))  severity failure;
	assert RAM(28709) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28709))))  severity failure;
	assert RAM(28710) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(28710))))  severity failure;
	assert RAM(28711) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(28711))))  severity failure;
	assert RAM(28712) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28712))))  severity failure;
	assert RAM(28713) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(28713))))  severity failure;
	assert RAM(28714) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28714))))  severity failure;
	assert RAM(28715) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28715))))  severity failure;
	assert RAM(28716) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28716))))  severity failure;
	assert RAM(28717) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(28717))))  severity failure;
	assert RAM(28718) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28718))))  severity failure;
	assert RAM(28719) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(28719))))  severity failure;
	assert RAM(28720) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28720))))  severity failure;
	assert RAM(28721) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(28721))))  severity failure;
	assert RAM(28722) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(28722))))  severity failure;
	assert RAM(28723) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28723))))  severity failure;
	assert RAM(28724) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28724))))  severity failure;
	assert RAM(28725) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(28725))))  severity failure;
	assert RAM(28726) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(28726))))  severity failure;
	assert RAM(28727) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(28727))))  severity failure;
	assert RAM(28728) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(28728))))  severity failure;
	assert RAM(28729) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(28729))))  severity failure;
	assert RAM(28730) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28730))))  severity failure;
	assert RAM(28731) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(28731))))  severity failure;
	assert RAM(28732) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28732))))  severity failure;
	assert RAM(28733) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28733))))  severity failure;
	assert RAM(28734) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(28734))))  severity failure;
	assert RAM(28735) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(28735))))  severity failure;
	assert RAM(28736) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(28736))))  severity failure;
	assert RAM(28737) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(28737))))  severity failure;
	assert RAM(28738) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(28738))))  severity failure;
	assert RAM(28739) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28739))))  severity failure;
	assert RAM(28740) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(28740))))  severity failure;
	assert RAM(28741) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(28741))))  severity failure;
	assert RAM(28742) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(28742))))  severity failure;
	assert RAM(28743) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(28743))))  severity failure;
	assert RAM(28744) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28744))))  severity failure;
	assert RAM(28745) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(28745))))  severity failure;
	assert RAM(28746) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28746))))  severity failure;
	assert RAM(28747) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(28747))))  severity failure;
	assert RAM(28748) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28748))))  severity failure;
	assert RAM(28749) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28749))))  severity failure;
	assert RAM(28750) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(28750))))  severity failure;
	assert RAM(28751) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(28751))))  severity failure;
	assert RAM(28752) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(28752))))  severity failure;
	assert RAM(28753) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(28753))))  severity failure;
	assert RAM(28754) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(28754))))  severity failure;
	assert RAM(28755) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(28755))))  severity failure;
	assert RAM(28756) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(28756))))  severity failure;
	assert RAM(28757) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28757))))  severity failure;
	assert RAM(28758) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28758))))  severity failure;
	assert RAM(28759) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(28759))))  severity failure;
	assert RAM(28760) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(28760))))  severity failure;
	assert RAM(28761) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(28761))))  severity failure;
	assert RAM(28762) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28762))))  severity failure;
	assert RAM(28763) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(28763))))  severity failure;
	assert RAM(28764) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(28764))))  severity failure;
	assert RAM(28765) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(28765))))  severity failure;
	assert RAM(28766) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(28766))))  severity failure;
	assert RAM(28767) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(28767))))  severity failure;
	assert RAM(28768) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28768))))  severity failure;
	assert RAM(28769) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28769))))  severity failure;
	assert RAM(28770) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(28770))))  severity failure;
	assert RAM(28771) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(28771))))  severity failure;
	assert RAM(28772) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28772))))  severity failure;
	assert RAM(28773) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(28773))))  severity failure;
	assert RAM(28774) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(28774))))  severity failure;
	assert RAM(28775) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(28775))))  severity failure;
	assert RAM(28776) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(28776))))  severity failure;
	assert RAM(28777) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(28777))))  severity failure;
	assert RAM(28778) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(28778))))  severity failure;
	assert RAM(28779) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(28779))))  severity failure;
	assert RAM(28780) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(28780))))  severity failure;
	assert RAM(28781) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(28781))))  severity failure;
	assert RAM(28782) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28782))))  severity failure;
	assert RAM(28783) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(28783))))  severity failure;
	assert RAM(28784) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28784))))  severity failure;
	assert RAM(28785) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28785))))  severity failure;
	assert RAM(28786) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(28786))))  severity failure;
	assert RAM(28787) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(28787))))  severity failure;
	assert RAM(28788) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(28788))))  severity failure;
	assert RAM(28789) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(28789))))  severity failure;
	assert RAM(28790) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(28790))))  severity failure;
	assert RAM(28791) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(28791))))  severity failure;
	assert RAM(28792) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28792))))  severity failure;
	assert RAM(28793) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(28793))))  severity failure;
	assert RAM(28794) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(28794))))  severity failure;
	assert RAM(28795) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28795))))  severity failure;
	assert RAM(28796) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28796))))  severity failure;
	assert RAM(28797) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(28797))))  severity failure;
	assert RAM(28798) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(28798))))  severity failure;
	assert RAM(28799) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(28799))))  severity failure;
	assert RAM(28800) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(28800))))  severity failure;
	assert RAM(28801) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(28801))))  severity failure;
	assert RAM(28802) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(28802))))  severity failure;
	assert RAM(28803) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(28803))))  severity failure;
	assert RAM(28804) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(28804))))  severity failure;
	assert RAM(28805) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(28805))))  severity failure;
	assert RAM(28806) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(28806))))  severity failure;
	assert RAM(28807) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28807))))  severity failure;
	assert RAM(28808) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(28808))))  severity failure;
	assert RAM(28809) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(28809))))  severity failure;
	assert RAM(28810) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(28810))))  severity failure;
	assert RAM(28811) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(28811))))  severity failure;
	assert RAM(28812) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(28812))))  severity failure;
	assert RAM(28813) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(28813))))  severity failure;
	assert RAM(28814) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(28814))))  severity failure;
	assert RAM(28815) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(28815))))  severity failure;
	assert RAM(28816) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(28816))))  severity failure;
	assert RAM(28817) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(28817))))  severity failure;
	assert RAM(28818) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(28818))))  severity failure;
	assert RAM(28819) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28819))))  severity failure;
	assert RAM(28820) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(28820))))  severity failure;
	assert RAM(28821) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(28821))))  severity failure;
	assert RAM(28822) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28822))))  severity failure;
	assert RAM(28823) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(28823))))  severity failure;
	assert RAM(28824) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28824))))  severity failure;
	assert RAM(28825) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(28825))))  severity failure;
	assert RAM(28826) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(28826))))  severity failure;
	assert RAM(28827) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28827))))  severity failure;
	assert RAM(28828) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28828))))  severity failure;
	assert RAM(28829) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28829))))  severity failure;
	assert RAM(28830) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(28830))))  severity failure;
	assert RAM(28831) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28831))))  severity failure;
	assert RAM(28832) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(28832))))  severity failure;
	assert RAM(28833) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(28833))))  severity failure;
	assert RAM(28834) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(28834))))  severity failure;
	assert RAM(28835) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28835))))  severity failure;
	assert RAM(28836) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(28836))))  severity failure;
	assert RAM(28837) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(28837))))  severity failure;
	assert RAM(28838) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28838))))  severity failure;
	assert RAM(28839) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(28839))))  severity failure;
	assert RAM(28840) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(28840))))  severity failure;
	assert RAM(28841) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(28841))))  severity failure;
	assert RAM(28842) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28842))))  severity failure;
	assert RAM(28843) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(28843))))  severity failure;
	assert RAM(28844) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(28844))))  severity failure;
	assert RAM(28845) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(28845))))  severity failure;
	assert RAM(28846) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(28846))))  severity failure;
	assert RAM(28847) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(28847))))  severity failure;
	assert RAM(28848) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28848))))  severity failure;
	assert RAM(28849) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(28849))))  severity failure;
	assert RAM(28850) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(28850))))  severity failure;
	assert RAM(28851) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28851))))  severity failure;
	assert RAM(28852) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(28852))))  severity failure;
	assert RAM(28853) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(28853))))  severity failure;
	assert RAM(28854) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(28854))))  severity failure;
	assert RAM(28855) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(28855))))  severity failure;
	assert RAM(28856) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(28856))))  severity failure;
	assert RAM(28857) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(28857))))  severity failure;
	assert RAM(28858) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(28858))))  severity failure;
	assert RAM(28859) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(28859))))  severity failure;
	assert RAM(28860) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28860))))  severity failure;
	assert RAM(28861) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(28861))))  severity failure;
	assert RAM(28862) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(28862))))  severity failure;
	assert RAM(28863) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(28863))))  severity failure;
	assert RAM(28864) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(28864))))  severity failure;
	assert RAM(28865) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28865))))  severity failure;
	assert RAM(28866) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(28866))))  severity failure;
	assert RAM(28867) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(28867))))  severity failure;
	assert RAM(28868) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(28868))))  severity failure;
	assert RAM(28869) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(28869))))  severity failure;
	assert RAM(28870) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(28870))))  severity failure;
	assert RAM(28871) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(28871))))  severity failure;
	assert RAM(28872) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(28872))))  severity failure;
	assert RAM(28873) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(28873))))  severity failure;
	assert RAM(28874) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(28874))))  severity failure;
	assert RAM(28875) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28875))))  severity failure;
	assert RAM(28876) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28876))))  severity failure;
	assert RAM(28877) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(28877))))  severity failure;
	assert RAM(28878) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(28878))))  severity failure;
	assert RAM(28879) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(28879))))  severity failure;
	assert RAM(28880) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(28880))))  severity failure;
	assert RAM(28881) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(28881))))  severity failure;
	assert RAM(28882) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(28882))))  severity failure;
	assert RAM(28883) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28883))))  severity failure;
	assert RAM(28884) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(28884))))  severity failure;
	assert RAM(28885) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28885))))  severity failure;
	assert RAM(28886) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28886))))  severity failure;
	assert RAM(28887) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(28887))))  severity failure;
	assert RAM(28888) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(28888))))  severity failure;
	assert RAM(28889) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(28889))))  severity failure;
	assert RAM(28890) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28890))))  severity failure;
	assert RAM(28891) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(28891))))  severity failure;
	assert RAM(28892) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(28892))))  severity failure;
	assert RAM(28893) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28893))))  severity failure;
	assert RAM(28894) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(28894))))  severity failure;
	assert RAM(28895) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(28895))))  severity failure;
	assert RAM(28896) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(28896))))  severity failure;
	assert RAM(28897) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(28897))))  severity failure;
	assert RAM(28898) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(28898))))  severity failure;
	assert RAM(28899) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(28899))))  severity failure;
	assert RAM(28900) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(28900))))  severity failure;
	assert RAM(28901) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(28901))))  severity failure;
	assert RAM(28902) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(28902))))  severity failure;
	assert RAM(28903) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(28903))))  severity failure;
	assert RAM(28904) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(28904))))  severity failure;
	assert RAM(28905) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28905))))  severity failure;
	assert RAM(28906) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(28906))))  severity failure;
	assert RAM(28907) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(28907))))  severity failure;
	assert RAM(28908) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(28908))))  severity failure;
	assert RAM(28909) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(28909))))  severity failure;
	assert RAM(28910) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(28910))))  severity failure;
	assert RAM(28911) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(28911))))  severity failure;
	assert RAM(28912) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(28912))))  severity failure;
	assert RAM(28913) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(28913))))  severity failure;
	assert RAM(28914) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(28914))))  severity failure;
	assert RAM(28915) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(28915))))  severity failure;
	assert RAM(28916) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(28916))))  severity failure;
	assert RAM(28917) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(28917))))  severity failure;
	assert RAM(28918) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(28918))))  severity failure;
	assert RAM(28919) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28919))))  severity failure;
	assert RAM(28920) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(28920))))  severity failure;
	assert RAM(28921) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28921))))  severity failure;
	assert RAM(28922) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(28922))))  severity failure;
	assert RAM(28923) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(28923))))  severity failure;
	assert RAM(28924) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28924))))  severity failure;
	assert RAM(28925) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(28925))))  severity failure;
	assert RAM(28926) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(28926))))  severity failure;
	assert RAM(28927) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(28927))))  severity failure;
	assert RAM(28928) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28928))))  severity failure;
	assert RAM(28929) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(28929))))  severity failure;
	assert RAM(28930) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(28930))))  severity failure;
	assert RAM(28931) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(28931))))  severity failure;
	assert RAM(28932) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(28932))))  severity failure;
	assert RAM(28933) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(28933))))  severity failure;
	assert RAM(28934) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(28934))))  severity failure;
	assert RAM(28935) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(28935))))  severity failure;
	assert RAM(28936) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(28936))))  severity failure;
	assert RAM(28937) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(28937))))  severity failure;
	assert RAM(28938) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(28938))))  severity failure;
	assert RAM(28939) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(28939))))  severity failure;
	assert RAM(28940) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(28940))))  severity failure;
	assert RAM(28941) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(28941))))  severity failure;
	assert RAM(28942) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(28942))))  severity failure;
	assert RAM(28943) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(28943))))  severity failure;
	assert RAM(28944) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(28944))))  severity failure;
	assert RAM(28945) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(28945))))  severity failure;
	assert RAM(28946) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(28946))))  severity failure;
	assert RAM(28947) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(28947))))  severity failure;
	assert RAM(28948) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(28948))))  severity failure;
	assert RAM(28949) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(28949))))  severity failure;
	assert RAM(28950) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(28950))))  severity failure;
	assert RAM(28951) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(28951))))  severity failure;
	assert RAM(28952) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(28952))))  severity failure;
	assert RAM(28953) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(28953))))  severity failure;
	assert RAM(28954) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(28954))))  severity failure;
	assert RAM(28955) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(28955))))  severity failure;
	assert RAM(28956) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(28956))))  severity failure;
	assert RAM(28957) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(28957))))  severity failure;
	assert RAM(28958) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(28958))))  severity failure;
	assert RAM(28959) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(28959))))  severity failure;
	assert RAM(28960) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(28960))))  severity failure;
	assert RAM(28961) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(28961))))  severity failure;
	assert RAM(28962) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28962))))  severity failure;
	assert RAM(28963) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(28963))))  severity failure;
	assert RAM(28964) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28964))))  severity failure;
	assert RAM(28965) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(28965))))  severity failure;
	assert RAM(28966) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(28966))))  severity failure;
	assert RAM(28967) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(28967))))  severity failure;
	assert RAM(28968) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(28968))))  severity failure;
	assert RAM(28969) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(28969))))  severity failure;
	assert RAM(28970) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(28970))))  severity failure;
	assert RAM(28971) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(28971))))  severity failure;
	assert RAM(28972) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(28972))))  severity failure;
	assert RAM(28973) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(28973))))  severity failure;
	assert RAM(28974) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(28974))))  severity failure;
	assert RAM(28975) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(28975))))  severity failure;
	assert RAM(28976) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(28976))))  severity failure;
	assert RAM(28977) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(28977))))  severity failure;
	assert RAM(28978) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(28978))))  severity failure;
	assert RAM(28979) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(28979))))  severity failure;
	assert RAM(28980) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(28980))))  severity failure;
	assert RAM(28981) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(28981))))  severity failure;
	assert RAM(28982) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(28982))))  severity failure;
	assert RAM(28983) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(28983))))  severity failure;
	assert RAM(28984) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(28984))))  severity failure;
	assert RAM(28985) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(28985))))  severity failure;
	assert RAM(28986) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(28986))))  severity failure;
	assert RAM(28987) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(28987))))  severity failure;
	assert RAM(28988) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(28988))))  severity failure;
	assert RAM(28989) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(28989))))  severity failure;
	assert RAM(28990) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(28990))))  severity failure;
	assert RAM(28991) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(28991))))  severity failure;
	assert RAM(28992) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(28992))))  severity failure;
	assert RAM(28993) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(28993))))  severity failure;
	assert RAM(28994) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(28994))))  severity failure;
	assert RAM(28995) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(28995))))  severity failure;
	assert RAM(28996) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(28996))))  severity failure;
	assert RAM(28997) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(28997))))  severity failure;
	assert RAM(28998) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(28998))))  severity failure;
	assert RAM(28999) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(28999))))  severity failure;
	assert RAM(29000) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(29000))))  severity failure;
	assert RAM(29001) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(29001))))  severity failure;
	assert RAM(29002) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29002))))  severity failure;
	assert RAM(29003) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29003))))  severity failure;
	assert RAM(29004) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(29004))))  severity failure;
	assert RAM(29005) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(29005))))  severity failure;
	assert RAM(29006) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29006))))  severity failure;
	assert RAM(29007) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29007))))  severity failure;
	assert RAM(29008) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(29008))))  severity failure;
	assert RAM(29009) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29009))))  severity failure;
	assert RAM(29010) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(29010))))  severity failure;
	assert RAM(29011) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29011))))  severity failure;
	assert RAM(29012) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29012))))  severity failure;
	assert RAM(29013) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29013))))  severity failure;
	assert RAM(29014) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(29014))))  severity failure;
	assert RAM(29015) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(29015))))  severity failure;
	assert RAM(29016) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29016))))  severity failure;
	assert RAM(29017) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(29017))))  severity failure;
	assert RAM(29018) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(29018))))  severity failure;
	assert RAM(29019) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(29019))))  severity failure;
	assert RAM(29020) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(29020))))  severity failure;
	assert RAM(29021) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(29021))))  severity failure;
	assert RAM(29022) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(29022))))  severity failure;
	assert RAM(29023) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(29023))))  severity failure;
	assert RAM(29024) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29024))))  severity failure;
	assert RAM(29025) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29025))))  severity failure;
	assert RAM(29026) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(29026))))  severity failure;
	assert RAM(29027) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(29027))))  severity failure;
	assert RAM(29028) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(29028))))  severity failure;
	assert RAM(29029) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29029))))  severity failure;
	assert RAM(29030) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29030))))  severity failure;
	assert RAM(29031) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29031))))  severity failure;
	assert RAM(29032) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(29032))))  severity failure;
	assert RAM(29033) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(29033))))  severity failure;
	assert RAM(29034) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(29034))))  severity failure;
	assert RAM(29035) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(29035))))  severity failure;
	assert RAM(29036) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29036))))  severity failure;
	assert RAM(29037) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29037))))  severity failure;
	assert RAM(29038) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(29038))))  severity failure;
	assert RAM(29039) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29039))))  severity failure;
	assert RAM(29040) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29040))))  severity failure;
	assert RAM(29041) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(29041))))  severity failure;
	assert RAM(29042) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(29042))))  severity failure;
	assert RAM(29043) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(29043))))  severity failure;
	assert RAM(29044) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(29044))))  severity failure;
	assert RAM(29045) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(29045))))  severity failure;
	assert RAM(29046) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(29046))))  severity failure;
	assert RAM(29047) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29047))))  severity failure;
	assert RAM(29048) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29048))))  severity failure;
	assert RAM(29049) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(29049))))  severity failure;
	assert RAM(29050) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(29050))))  severity failure;
	assert RAM(29051) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29051))))  severity failure;
	assert RAM(29052) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29052))))  severity failure;
	assert RAM(29053) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(29053))))  severity failure;
	assert RAM(29054) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(29054))))  severity failure;
	assert RAM(29055) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(29055))))  severity failure;
	assert RAM(29056) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(29056))))  severity failure;
	assert RAM(29057) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29057))))  severity failure;
	assert RAM(29058) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(29058))))  severity failure;
	assert RAM(29059) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(29059))))  severity failure;
	assert RAM(29060) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29060))))  severity failure;
	assert RAM(29061) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(29061))))  severity failure;
	assert RAM(29062) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(29062))))  severity failure;
	assert RAM(29063) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29063))))  severity failure;
	assert RAM(29064) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(29064))))  severity failure;
	assert RAM(29065) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(29065))))  severity failure;
	assert RAM(29066) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(29066))))  severity failure;
	assert RAM(29067) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(29067))))  severity failure;
	assert RAM(29068) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(29068))))  severity failure;
	assert RAM(29069) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(29069))))  severity failure;
	assert RAM(29070) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29070))))  severity failure;
	assert RAM(29071) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(29071))))  severity failure;
	assert RAM(29072) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29072))))  severity failure;
	assert RAM(29073) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(29073))))  severity failure;
	assert RAM(29074) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(29074))))  severity failure;
	assert RAM(29075) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29075))))  severity failure;
	assert RAM(29076) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29076))))  severity failure;
	assert RAM(29077) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29077))))  severity failure;
	assert RAM(29078) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29078))))  severity failure;
	assert RAM(29079) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(29079))))  severity failure;
	assert RAM(29080) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29080))))  severity failure;
	assert RAM(29081) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(29081))))  severity failure;
	assert RAM(29082) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29082))))  severity failure;
	assert RAM(29083) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29083))))  severity failure;
	assert RAM(29084) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29084))))  severity failure;
	assert RAM(29085) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(29085))))  severity failure;
	assert RAM(29086) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(29086))))  severity failure;
	assert RAM(29087) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(29087))))  severity failure;
	assert RAM(29088) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29088))))  severity failure;
	assert RAM(29089) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(29089))))  severity failure;
	assert RAM(29090) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29090))))  severity failure;
	assert RAM(29091) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(29091))))  severity failure;
	assert RAM(29092) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(29092))))  severity failure;
	assert RAM(29093) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29093))))  severity failure;
	assert RAM(29094) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(29094))))  severity failure;
	assert RAM(29095) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(29095))))  severity failure;
	assert RAM(29096) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(29096))))  severity failure;
	assert RAM(29097) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29097))))  severity failure;
	assert RAM(29098) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(29098))))  severity failure;
	assert RAM(29099) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(29099))))  severity failure;
	assert RAM(29100) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(29100))))  severity failure;
	assert RAM(29101) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29101))))  severity failure;
	assert RAM(29102) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29102))))  severity failure;
	assert RAM(29103) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(29103))))  severity failure;
	assert RAM(29104) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(29104))))  severity failure;
	assert RAM(29105) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(29105))))  severity failure;
	assert RAM(29106) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29106))))  severity failure;
	assert RAM(29107) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29107))))  severity failure;
	assert RAM(29108) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29108))))  severity failure;
	assert RAM(29109) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29109))))  severity failure;
	assert RAM(29110) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(29110))))  severity failure;
	assert RAM(29111) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(29111))))  severity failure;
	assert RAM(29112) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29112))))  severity failure;
	assert RAM(29113) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(29113))))  severity failure;
	assert RAM(29114) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(29114))))  severity failure;
	assert RAM(29115) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(29115))))  severity failure;
	assert RAM(29116) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29116))))  severity failure;
	assert RAM(29117) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(29117))))  severity failure;
	assert RAM(29118) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(29118))))  severity failure;
	assert RAM(29119) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(29119))))  severity failure;
	assert RAM(29120) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(29120))))  severity failure;
	assert RAM(29121) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(29121))))  severity failure;
	assert RAM(29122) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(29122))))  severity failure;
	assert RAM(29123) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(29123))))  severity failure;
	assert RAM(29124) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(29124))))  severity failure;
	assert RAM(29125) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(29125))))  severity failure;
	assert RAM(29126) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(29126))))  severity failure;
	assert RAM(29127) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29127))))  severity failure;
	assert RAM(29128) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(29128))))  severity failure;
	assert RAM(29129) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(29129))))  severity failure;
	assert RAM(29130) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(29130))))  severity failure;
	assert RAM(29131) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(29131))))  severity failure;
	assert RAM(29132) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29132))))  severity failure;
	assert RAM(29133) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(29133))))  severity failure;
	assert RAM(29134) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(29134))))  severity failure;
	assert RAM(29135) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29135))))  severity failure;
	assert RAM(29136) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(29136))))  severity failure;
	assert RAM(29137) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(29137))))  severity failure;
	assert RAM(29138) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(29138))))  severity failure;
	assert RAM(29139) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29139))))  severity failure;
	assert RAM(29140) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(29140))))  severity failure;
	assert RAM(29141) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(29141))))  severity failure;
	assert RAM(29142) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29142))))  severity failure;
	assert RAM(29143) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(29143))))  severity failure;
	assert RAM(29144) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(29144))))  severity failure;
	assert RAM(29145) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(29145))))  severity failure;
	assert RAM(29146) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(29146))))  severity failure;
	assert RAM(29147) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(29147))))  severity failure;
	assert RAM(29148) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(29148))))  severity failure;
	assert RAM(29149) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29149))))  severity failure;
	assert RAM(29150) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29150))))  severity failure;
	assert RAM(29151) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(29151))))  severity failure;
	assert RAM(29152) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(29152))))  severity failure;
	assert RAM(29153) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(29153))))  severity failure;
	assert RAM(29154) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(29154))))  severity failure;
	assert RAM(29155) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29155))))  severity failure;
	assert RAM(29156) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29156))))  severity failure;
	assert RAM(29157) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29157))))  severity failure;
	assert RAM(29158) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(29158))))  severity failure;
	assert RAM(29159) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(29159))))  severity failure;
	assert RAM(29160) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(29160))))  severity failure;
	assert RAM(29161) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(29161))))  severity failure;
	assert RAM(29162) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(29162))))  severity failure;
	assert RAM(29163) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(29163))))  severity failure;
	assert RAM(29164) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(29164))))  severity failure;
	assert RAM(29165) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(29165))))  severity failure;
	assert RAM(29166) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29166))))  severity failure;
	assert RAM(29167) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(29167))))  severity failure;
	assert RAM(29168) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(29168))))  severity failure;
	assert RAM(29169) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(29169))))  severity failure;
	assert RAM(29170) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29170))))  severity failure;
	assert RAM(29171) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29171))))  severity failure;
	assert RAM(29172) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29172))))  severity failure;
	assert RAM(29173) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(29173))))  severity failure;
	assert RAM(29174) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29174))))  severity failure;
	assert RAM(29175) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(29175))))  severity failure;
	assert RAM(29176) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(29176))))  severity failure;
	assert RAM(29177) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(29177))))  severity failure;
	assert RAM(29178) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(29178))))  severity failure;
	assert RAM(29179) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29179))))  severity failure;
	assert RAM(29180) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(29180))))  severity failure;
	assert RAM(29181) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(29181))))  severity failure;
	assert RAM(29182) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(29182))))  severity failure;
	assert RAM(29183) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29183))))  severity failure;
	assert RAM(29184) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(29184))))  severity failure;
	assert RAM(29185) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(29185))))  severity failure;
	assert RAM(29186) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29186))))  severity failure;
	assert RAM(29187) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29187))))  severity failure;
	assert RAM(29188) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(29188))))  severity failure;
	assert RAM(29189) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29189))))  severity failure;
	assert RAM(29190) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(29190))))  severity failure;
	assert RAM(29191) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(29191))))  severity failure;
	assert RAM(29192) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(29192))))  severity failure;
	assert RAM(29193) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(29193))))  severity failure;
	assert RAM(29194) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(29194))))  severity failure;
	assert RAM(29195) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(29195))))  severity failure;
	assert RAM(29196) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29196))))  severity failure;
	assert RAM(29197) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(29197))))  severity failure;
	assert RAM(29198) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29198))))  severity failure;
	assert RAM(29199) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(29199))))  severity failure;
	assert RAM(29200) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29200))))  severity failure;
	assert RAM(29201) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29201))))  severity failure;
	assert RAM(29202) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29202))))  severity failure;
	assert RAM(29203) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(29203))))  severity failure;
	assert RAM(29204) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(29204))))  severity failure;
	assert RAM(29205) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(29205))))  severity failure;
	assert RAM(29206) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29206))))  severity failure;
	assert RAM(29207) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(29207))))  severity failure;
	assert RAM(29208) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(29208))))  severity failure;
	assert RAM(29209) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(29209))))  severity failure;
	assert RAM(29210) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(29210))))  severity failure;
	assert RAM(29211) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(29211))))  severity failure;
	assert RAM(29212) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(29212))))  severity failure;
	assert RAM(29213) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(29213))))  severity failure;
	assert RAM(29214) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(29214))))  severity failure;
	assert RAM(29215) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29215))))  severity failure;
	assert RAM(29216) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(29216))))  severity failure;
	assert RAM(29217) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29217))))  severity failure;
	assert RAM(29218) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(29218))))  severity failure;
	assert RAM(29219) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(29219))))  severity failure;
	assert RAM(29220) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(29220))))  severity failure;
	assert RAM(29221) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29221))))  severity failure;
	assert RAM(29222) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29222))))  severity failure;
	assert RAM(29223) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29223))))  severity failure;
	assert RAM(29224) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(29224))))  severity failure;
	assert RAM(29225) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(29225))))  severity failure;
	assert RAM(29226) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(29226))))  severity failure;
	assert RAM(29227) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(29227))))  severity failure;
	assert RAM(29228) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29228))))  severity failure;
	assert RAM(29229) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29229))))  severity failure;
	assert RAM(29230) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29230))))  severity failure;
	assert RAM(29231) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29231))))  severity failure;
	assert RAM(29232) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(29232))))  severity failure;
	assert RAM(29233) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(29233))))  severity failure;
	assert RAM(29234) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(29234))))  severity failure;
	assert RAM(29235) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(29235))))  severity failure;
	assert RAM(29236) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(29236))))  severity failure;
	assert RAM(29237) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(29237))))  severity failure;
	assert RAM(29238) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(29238))))  severity failure;
	assert RAM(29239) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29239))))  severity failure;
	assert RAM(29240) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(29240))))  severity failure;
	assert RAM(29241) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(29241))))  severity failure;
	assert RAM(29242) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29242))))  severity failure;
	assert RAM(29243) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(29243))))  severity failure;
	assert RAM(29244) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29244))))  severity failure;
	assert RAM(29245) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29245))))  severity failure;
	assert RAM(29246) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(29246))))  severity failure;
	assert RAM(29247) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(29247))))  severity failure;
	assert RAM(29248) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29248))))  severity failure;
	assert RAM(29249) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(29249))))  severity failure;
	assert RAM(29250) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29250))))  severity failure;
	assert RAM(29251) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(29251))))  severity failure;
	assert RAM(29252) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(29252))))  severity failure;
	assert RAM(29253) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29253))))  severity failure;
	assert RAM(29254) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29254))))  severity failure;
	assert RAM(29255) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29255))))  severity failure;
	assert RAM(29256) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29256))))  severity failure;
	assert RAM(29257) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29257))))  severity failure;
	assert RAM(29258) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29258))))  severity failure;
	assert RAM(29259) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29259))))  severity failure;
	assert RAM(29260) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(29260))))  severity failure;
	assert RAM(29261) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(29261))))  severity failure;
	assert RAM(29262) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(29262))))  severity failure;
	assert RAM(29263) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29263))))  severity failure;
	assert RAM(29264) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29264))))  severity failure;
	assert RAM(29265) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29265))))  severity failure;
	assert RAM(29266) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29266))))  severity failure;
	assert RAM(29267) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(29267))))  severity failure;
	assert RAM(29268) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(29268))))  severity failure;
	assert RAM(29269) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(29269))))  severity failure;
	assert RAM(29270) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29270))))  severity failure;
	assert RAM(29271) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29271))))  severity failure;
	assert RAM(29272) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29272))))  severity failure;
	assert RAM(29273) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(29273))))  severity failure;
	assert RAM(29274) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(29274))))  severity failure;
	assert RAM(29275) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29275))))  severity failure;
	assert RAM(29276) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29276))))  severity failure;
	assert RAM(29277) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(29277))))  severity failure;
	assert RAM(29278) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(29278))))  severity failure;
	assert RAM(29279) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29279))))  severity failure;
	assert RAM(29280) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(29280))))  severity failure;
	assert RAM(29281) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29281))))  severity failure;
	assert RAM(29282) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(29282))))  severity failure;
	assert RAM(29283) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29283))))  severity failure;
	assert RAM(29284) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(29284))))  severity failure;
	assert RAM(29285) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29285))))  severity failure;
	assert RAM(29286) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(29286))))  severity failure;
	assert RAM(29287) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(29287))))  severity failure;
	assert RAM(29288) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(29288))))  severity failure;
	assert RAM(29289) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(29289))))  severity failure;
	assert RAM(29290) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(29290))))  severity failure;
	assert RAM(29291) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29291))))  severity failure;
	assert RAM(29292) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29292))))  severity failure;
	assert RAM(29293) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29293))))  severity failure;
	assert RAM(29294) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29294))))  severity failure;
	assert RAM(29295) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(29295))))  severity failure;
	assert RAM(29296) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(29296))))  severity failure;
	assert RAM(29297) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(29297))))  severity failure;
	assert RAM(29298) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29298))))  severity failure;
	assert RAM(29299) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(29299))))  severity failure;
	assert RAM(29300) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(29300))))  severity failure;
	assert RAM(29301) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(29301))))  severity failure;
	assert RAM(29302) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(29302))))  severity failure;
	assert RAM(29303) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(29303))))  severity failure;
	assert RAM(29304) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(29304))))  severity failure;
	assert RAM(29305) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(29305))))  severity failure;
	assert RAM(29306) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(29306))))  severity failure;
	assert RAM(29307) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29307))))  severity failure;
	assert RAM(29308) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(29308))))  severity failure;
	assert RAM(29309) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(29309))))  severity failure;
	assert RAM(29310) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29310))))  severity failure;
	assert RAM(29311) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29311))))  severity failure;
	assert RAM(29312) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29312))))  severity failure;
	assert RAM(29313) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29313))))  severity failure;
	assert RAM(29314) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29314))))  severity failure;
	assert RAM(29315) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(29315))))  severity failure;
	assert RAM(29316) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(29316))))  severity failure;
	assert RAM(29317) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(29317))))  severity failure;
	assert RAM(29318) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(29318))))  severity failure;
	assert RAM(29319) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29319))))  severity failure;
	assert RAM(29320) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29320))))  severity failure;
	assert RAM(29321) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29321))))  severity failure;
	assert RAM(29322) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(29322))))  severity failure;
	assert RAM(29323) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(29323))))  severity failure;
	assert RAM(29324) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29324))))  severity failure;
	assert RAM(29325) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(29325))))  severity failure;
	assert RAM(29326) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(29326))))  severity failure;
	assert RAM(29327) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(29327))))  severity failure;
	assert RAM(29328) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29328))))  severity failure;
	assert RAM(29329) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(29329))))  severity failure;
	assert RAM(29330) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(29330))))  severity failure;
	assert RAM(29331) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29331))))  severity failure;
	assert RAM(29332) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29332))))  severity failure;
	assert RAM(29333) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29333))))  severity failure;
	assert RAM(29334) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29334))))  severity failure;
	assert RAM(29335) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(29335))))  severity failure;
	assert RAM(29336) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(29336))))  severity failure;
	assert RAM(29337) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(29337))))  severity failure;
	assert RAM(29338) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(29338))))  severity failure;
	assert RAM(29339) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(29339))))  severity failure;
	assert RAM(29340) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(29340))))  severity failure;
	assert RAM(29341) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(29341))))  severity failure;
	assert RAM(29342) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(29342))))  severity failure;
	assert RAM(29343) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29343))))  severity failure;
	assert RAM(29344) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(29344))))  severity failure;
	assert RAM(29345) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(29345))))  severity failure;
	assert RAM(29346) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(29346))))  severity failure;
	assert RAM(29347) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(29347))))  severity failure;
	assert RAM(29348) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29348))))  severity failure;
	assert RAM(29349) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29349))))  severity failure;
	assert RAM(29350) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(29350))))  severity failure;
	assert RAM(29351) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(29351))))  severity failure;
	assert RAM(29352) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29352))))  severity failure;
	assert RAM(29353) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29353))))  severity failure;
	assert RAM(29354) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(29354))))  severity failure;
	assert RAM(29355) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(29355))))  severity failure;
	assert RAM(29356) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29356))))  severity failure;
	assert RAM(29357) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(29357))))  severity failure;
	assert RAM(29358) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(29358))))  severity failure;
	assert RAM(29359) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29359))))  severity failure;
	assert RAM(29360) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(29360))))  severity failure;
	assert RAM(29361) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(29361))))  severity failure;
	assert RAM(29362) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(29362))))  severity failure;
	assert RAM(29363) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(29363))))  severity failure;
	assert RAM(29364) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(29364))))  severity failure;
	assert RAM(29365) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(29365))))  severity failure;
	assert RAM(29366) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29366))))  severity failure;
	assert RAM(29367) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(29367))))  severity failure;
	assert RAM(29368) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(29368))))  severity failure;
	assert RAM(29369) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29369))))  severity failure;
	assert RAM(29370) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29370))))  severity failure;
	assert RAM(29371) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29371))))  severity failure;
	assert RAM(29372) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(29372))))  severity failure;
	assert RAM(29373) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29373))))  severity failure;
	assert RAM(29374) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(29374))))  severity failure;
	assert RAM(29375) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(29375))))  severity failure;
	assert RAM(29376) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(29376))))  severity failure;
	assert RAM(29377) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(29377))))  severity failure;
	assert RAM(29378) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(29378))))  severity failure;
	assert RAM(29379) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(29379))))  severity failure;
	assert RAM(29380) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(29380))))  severity failure;
	assert RAM(29381) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(29381))))  severity failure;
	assert RAM(29382) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29382))))  severity failure;
	assert RAM(29383) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(29383))))  severity failure;
	assert RAM(29384) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(29384))))  severity failure;
	assert RAM(29385) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(29385))))  severity failure;
	assert RAM(29386) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29386))))  severity failure;
	assert RAM(29387) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29387))))  severity failure;
	assert RAM(29388) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29388))))  severity failure;
	assert RAM(29389) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(29389))))  severity failure;
	assert RAM(29390) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29390))))  severity failure;
	assert RAM(29391) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(29391))))  severity failure;
	assert RAM(29392) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(29392))))  severity failure;
	assert RAM(29393) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29393))))  severity failure;
	assert RAM(29394) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29394))))  severity failure;
	assert RAM(29395) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(29395))))  severity failure;
	assert RAM(29396) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(29396))))  severity failure;
	assert RAM(29397) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(29397))))  severity failure;
	assert RAM(29398) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29398))))  severity failure;
	assert RAM(29399) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(29399))))  severity failure;
	assert RAM(29400) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(29400))))  severity failure;
	assert RAM(29401) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29401))))  severity failure;
	assert RAM(29402) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(29402))))  severity failure;
	assert RAM(29403) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(29403))))  severity failure;
	assert RAM(29404) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29404))))  severity failure;
	assert RAM(29405) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29405))))  severity failure;
	assert RAM(29406) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(29406))))  severity failure;
	assert RAM(29407) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29407))))  severity failure;
	assert RAM(29408) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29408))))  severity failure;
	assert RAM(29409) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(29409))))  severity failure;
	assert RAM(29410) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(29410))))  severity failure;
	assert RAM(29411) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(29411))))  severity failure;
	assert RAM(29412) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(29412))))  severity failure;
	assert RAM(29413) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(29413))))  severity failure;
	assert RAM(29414) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29414))))  severity failure;
	assert RAM(29415) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(29415))))  severity failure;
	assert RAM(29416) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(29416))))  severity failure;
	assert RAM(29417) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(29417))))  severity failure;
	assert RAM(29418) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(29418))))  severity failure;
	assert RAM(29419) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(29419))))  severity failure;
	assert RAM(29420) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29420))))  severity failure;
	assert RAM(29421) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(29421))))  severity failure;
	assert RAM(29422) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29422))))  severity failure;
	assert RAM(29423) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(29423))))  severity failure;
	assert RAM(29424) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(29424))))  severity failure;
	assert RAM(29425) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(29425))))  severity failure;
	assert RAM(29426) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(29426))))  severity failure;
	assert RAM(29427) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29427))))  severity failure;
	assert RAM(29428) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(29428))))  severity failure;
	assert RAM(29429) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29429))))  severity failure;
	assert RAM(29430) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(29430))))  severity failure;
	assert RAM(29431) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29431))))  severity failure;
	assert RAM(29432) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(29432))))  severity failure;
	assert RAM(29433) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(29433))))  severity failure;
	assert RAM(29434) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(29434))))  severity failure;
	assert RAM(29435) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(29435))))  severity failure;
	assert RAM(29436) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(29436))))  severity failure;
	assert RAM(29437) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(29437))))  severity failure;
	assert RAM(29438) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29438))))  severity failure;
	assert RAM(29439) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(29439))))  severity failure;
	assert RAM(29440) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(29440))))  severity failure;
	assert RAM(29441) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(29441))))  severity failure;
	assert RAM(29442) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(29442))))  severity failure;
	assert RAM(29443) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(29443))))  severity failure;
	assert RAM(29444) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29444))))  severity failure;
	assert RAM(29445) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29445))))  severity failure;
	assert RAM(29446) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29446))))  severity failure;
	assert RAM(29447) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(29447))))  severity failure;
	assert RAM(29448) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(29448))))  severity failure;
	assert RAM(29449) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(29449))))  severity failure;
	assert RAM(29450) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29450))))  severity failure;
	assert RAM(29451) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(29451))))  severity failure;
	assert RAM(29452) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29452))))  severity failure;
	assert RAM(29453) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(29453))))  severity failure;
	assert RAM(29454) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(29454))))  severity failure;
	assert RAM(29455) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(29455))))  severity failure;
	assert RAM(29456) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(29456))))  severity failure;
	assert RAM(29457) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29457))))  severity failure;
	assert RAM(29458) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29458))))  severity failure;
	assert RAM(29459) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(29459))))  severity failure;
	assert RAM(29460) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29460))))  severity failure;
	assert RAM(29461) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(29461))))  severity failure;
	assert RAM(29462) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(29462))))  severity failure;
	assert RAM(29463) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29463))))  severity failure;
	assert RAM(29464) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(29464))))  severity failure;
	assert RAM(29465) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(29465))))  severity failure;
	assert RAM(29466) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(29466))))  severity failure;
	assert RAM(29467) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(29467))))  severity failure;
	assert RAM(29468) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(29468))))  severity failure;
	assert RAM(29469) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(29469))))  severity failure;
	assert RAM(29470) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29470))))  severity failure;
	assert RAM(29471) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29471))))  severity failure;
	assert RAM(29472) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(29472))))  severity failure;
	assert RAM(29473) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29473))))  severity failure;
	assert RAM(29474) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29474))))  severity failure;
	assert RAM(29475) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29475))))  severity failure;
	assert RAM(29476) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29476))))  severity failure;
	assert RAM(29477) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29477))))  severity failure;
	assert RAM(29478) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(29478))))  severity failure;
	assert RAM(29479) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29479))))  severity failure;
	assert RAM(29480) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(29480))))  severity failure;
	assert RAM(29481) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29481))))  severity failure;
	assert RAM(29482) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29482))))  severity failure;
	assert RAM(29483) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(29483))))  severity failure;
	assert RAM(29484) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(29484))))  severity failure;
	assert RAM(29485) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29485))))  severity failure;
	assert RAM(29486) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29486))))  severity failure;
	assert RAM(29487) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(29487))))  severity failure;
	assert RAM(29488) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(29488))))  severity failure;
	assert RAM(29489) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29489))))  severity failure;
	assert RAM(29490) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(29490))))  severity failure;
	assert RAM(29491) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(29491))))  severity failure;
	assert RAM(29492) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(29492))))  severity failure;
	assert RAM(29493) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29493))))  severity failure;
	assert RAM(29494) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(29494))))  severity failure;
	assert RAM(29495) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29495))))  severity failure;
	assert RAM(29496) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(29496))))  severity failure;
	assert RAM(29497) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(29497))))  severity failure;
	assert RAM(29498) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29498))))  severity failure;
	assert RAM(29499) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29499))))  severity failure;
	assert RAM(29500) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(29500))))  severity failure;
	assert RAM(29501) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(29501))))  severity failure;
	assert RAM(29502) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(29502))))  severity failure;
	assert RAM(29503) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29503))))  severity failure;
	assert RAM(29504) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(29504))))  severity failure;
	assert RAM(29505) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(29505))))  severity failure;
	assert RAM(29506) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(29506))))  severity failure;
	assert RAM(29507) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29507))))  severity failure;
	assert RAM(29508) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(29508))))  severity failure;
	assert RAM(29509) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(29509))))  severity failure;
	assert RAM(29510) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(29510))))  severity failure;
	assert RAM(29511) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(29511))))  severity failure;
	assert RAM(29512) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(29512))))  severity failure;
	assert RAM(29513) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29513))))  severity failure;
	assert RAM(29514) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29514))))  severity failure;
	assert RAM(29515) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29515))))  severity failure;
	assert RAM(29516) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(29516))))  severity failure;
	assert RAM(29517) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(29517))))  severity failure;
	assert RAM(29518) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29518))))  severity failure;
	assert RAM(29519) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(29519))))  severity failure;
	assert RAM(29520) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29520))))  severity failure;
	assert RAM(29521) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(29521))))  severity failure;
	assert RAM(29522) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(29522))))  severity failure;
	assert RAM(29523) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(29523))))  severity failure;
	assert RAM(29524) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(29524))))  severity failure;
	assert RAM(29525) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(29525))))  severity failure;
	assert RAM(29526) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(29526))))  severity failure;
	assert RAM(29527) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29527))))  severity failure;
	assert RAM(29528) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(29528))))  severity failure;
	assert RAM(29529) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29529))))  severity failure;
	assert RAM(29530) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(29530))))  severity failure;
	assert RAM(29531) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29531))))  severity failure;
	assert RAM(29532) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(29532))))  severity failure;
	assert RAM(29533) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(29533))))  severity failure;
	assert RAM(29534) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29534))))  severity failure;
	assert RAM(29535) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(29535))))  severity failure;
	assert RAM(29536) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29536))))  severity failure;
	assert RAM(29537) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29537))))  severity failure;
	assert RAM(29538) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(29538))))  severity failure;
	assert RAM(29539) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29539))))  severity failure;
	assert RAM(29540) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29540))))  severity failure;
	assert RAM(29541) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29541))))  severity failure;
	assert RAM(29542) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(29542))))  severity failure;
	assert RAM(29543) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(29543))))  severity failure;
	assert RAM(29544) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(29544))))  severity failure;
	assert RAM(29545) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(29545))))  severity failure;
	assert RAM(29546) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(29546))))  severity failure;
	assert RAM(29547) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29547))))  severity failure;
	assert RAM(29548) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(29548))))  severity failure;
	assert RAM(29549) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(29549))))  severity failure;
	assert RAM(29550) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(29550))))  severity failure;
	assert RAM(29551) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(29551))))  severity failure;
	assert RAM(29552) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(29552))))  severity failure;
	assert RAM(29553) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29553))))  severity failure;
	assert RAM(29554) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(29554))))  severity failure;
	assert RAM(29555) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29555))))  severity failure;
	assert RAM(29556) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29556))))  severity failure;
	assert RAM(29557) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29557))))  severity failure;
	assert RAM(29558) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(29558))))  severity failure;
	assert RAM(29559) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(29559))))  severity failure;
	assert RAM(29560) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(29560))))  severity failure;
	assert RAM(29561) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29561))))  severity failure;
	assert RAM(29562) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(29562))))  severity failure;
	assert RAM(29563) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29563))))  severity failure;
	assert RAM(29564) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29564))))  severity failure;
	assert RAM(29565) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(29565))))  severity failure;
	assert RAM(29566) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(29566))))  severity failure;
	assert RAM(29567) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(29567))))  severity failure;
	assert RAM(29568) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29568))))  severity failure;
	assert RAM(29569) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(29569))))  severity failure;
	assert RAM(29570) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29570))))  severity failure;
	assert RAM(29571) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(29571))))  severity failure;
	assert RAM(29572) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(29572))))  severity failure;
	assert RAM(29573) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(29573))))  severity failure;
	assert RAM(29574) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(29574))))  severity failure;
	assert RAM(29575) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(29575))))  severity failure;
	assert RAM(29576) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29576))))  severity failure;
	assert RAM(29577) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29577))))  severity failure;
	assert RAM(29578) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29578))))  severity failure;
	assert RAM(29579) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29579))))  severity failure;
	assert RAM(29580) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29580))))  severity failure;
	assert RAM(29581) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29581))))  severity failure;
	assert RAM(29582) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(29582))))  severity failure;
	assert RAM(29583) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(29583))))  severity failure;
	assert RAM(29584) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(29584))))  severity failure;
	assert RAM(29585) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(29585))))  severity failure;
	assert RAM(29586) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29586))))  severity failure;
	assert RAM(29587) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(29587))))  severity failure;
	assert RAM(29588) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(29588))))  severity failure;
	assert RAM(29589) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(29589))))  severity failure;
	assert RAM(29590) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29590))))  severity failure;
	assert RAM(29591) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(29591))))  severity failure;
	assert RAM(29592) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29592))))  severity failure;
	assert RAM(29593) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(29593))))  severity failure;
	assert RAM(29594) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(29594))))  severity failure;
	assert RAM(29595) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29595))))  severity failure;
	assert RAM(29596) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29596))))  severity failure;
	assert RAM(29597) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(29597))))  severity failure;
	assert RAM(29598) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(29598))))  severity failure;
	assert RAM(29599) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(29599))))  severity failure;
	assert RAM(29600) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(29600))))  severity failure;
	assert RAM(29601) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(29601))))  severity failure;
	assert RAM(29602) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29602))))  severity failure;
	assert RAM(29603) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29603))))  severity failure;
	assert RAM(29604) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(29604))))  severity failure;
	assert RAM(29605) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(29605))))  severity failure;
	assert RAM(29606) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29606))))  severity failure;
	assert RAM(29607) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29607))))  severity failure;
	assert RAM(29608) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(29608))))  severity failure;
	assert RAM(29609) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(29609))))  severity failure;
	assert RAM(29610) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(29610))))  severity failure;
	assert RAM(29611) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(29611))))  severity failure;
	assert RAM(29612) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(29612))))  severity failure;
	assert RAM(29613) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29613))))  severity failure;
	assert RAM(29614) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(29614))))  severity failure;
	assert RAM(29615) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(29615))))  severity failure;
	assert RAM(29616) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(29616))))  severity failure;
	assert RAM(29617) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29617))))  severity failure;
	assert RAM(29618) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(29618))))  severity failure;
	assert RAM(29619) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(29619))))  severity failure;
	assert RAM(29620) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(29620))))  severity failure;
	assert RAM(29621) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29621))))  severity failure;
	assert RAM(29622) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29622))))  severity failure;
	assert RAM(29623) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(29623))))  severity failure;
	assert RAM(29624) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29624))))  severity failure;
	assert RAM(29625) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(29625))))  severity failure;
	assert RAM(29626) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(29626))))  severity failure;
	assert RAM(29627) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29627))))  severity failure;
	assert RAM(29628) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29628))))  severity failure;
	assert RAM(29629) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(29629))))  severity failure;
	assert RAM(29630) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(29630))))  severity failure;
	assert RAM(29631) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29631))))  severity failure;
	assert RAM(29632) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(29632))))  severity failure;
	assert RAM(29633) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29633))))  severity failure;
	assert RAM(29634) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(29634))))  severity failure;
	assert RAM(29635) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(29635))))  severity failure;
	assert RAM(29636) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29636))))  severity failure;
	assert RAM(29637) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(29637))))  severity failure;
	assert RAM(29638) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(29638))))  severity failure;
	assert RAM(29639) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(29639))))  severity failure;
	assert RAM(29640) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29640))))  severity failure;
	assert RAM(29641) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(29641))))  severity failure;
	assert RAM(29642) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(29642))))  severity failure;
	assert RAM(29643) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29643))))  severity failure;
	assert RAM(29644) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(29644))))  severity failure;
	assert RAM(29645) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29645))))  severity failure;
	assert RAM(29646) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29646))))  severity failure;
	assert RAM(29647) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29647))))  severity failure;
	assert RAM(29648) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(29648))))  severity failure;
	assert RAM(29649) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(29649))))  severity failure;
	assert RAM(29650) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29650))))  severity failure;
	assert RAM(29651) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(29651))))  severity failure;
	assert RAM(29652) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29652))))  severity failure;
	assert RAM(29653) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(29653))))  severity failure;
	assert RAM(29654) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29654))))  severity failure;
	assert RAM(29655) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(29655))))  severity failure;
	assert RAM(29656) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(29656))))  severity failure;
	assert RAM(29657) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(29657))))  severity failure;
	assert RAM(29658) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29658))))  severity failure;
	assert RAM(29659) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29659))))  severity failure;
	assert RAM(29660) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(29660))))  severity failure;
	assert RAM(29661) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(29661))))  severity failure;
	assert RAM(29662) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29662))))  severity failure;
	assert RAM(29663) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29663))))  severity failure;
	assert RAM(29664) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(29664))))  severity failure;
	assert RAM(29665) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(29665))))  severity failure;
	assert RAM(29666) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(29666))))  severity failure;
	assert RAM(29667) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(29667))))  severity failure;
	assert RAM(29668) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(29668))))  severity failure;
	assert RAM(29669) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29669))))  severity failure;
	assert RAM(29670) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(29670))))  severity failure;
	assert RAM(29671) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(29671))))  severity failure;
	assert RAM(29672) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29672))))  severity failure;
	assert RAM(29673) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(29673))))  severity failure;
	assert RAM(29674) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29674))))  severity failure;
	assert RAM(29675) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(29675))))  severity failure;
	assert RAM(29676) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(29676))))  severity failure;
	assert RAM(29677) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(29677))))  severity failure;
	assert RAM(29678) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29678))))  severity failure;
	assert RAM(29679) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29679))))  severity failure;
	assert RAM(29680) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(29680))))  severity failure;
	assert RAM(29681) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29681))))  severity failure;
	assert RAM(29682) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29682))))  severity failure;
	assert RAM(29683) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(29683))))  severity failure;
	assert RAM(29684) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(29684))))  severity failure;
	assert RAM(29685) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29685))))  severity failure;
	assert RAM(29686) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(29686))))  severity failure;
	assert RAM(29687) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(29687))))  severity failure;
	assert RAM(29688) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(29688))))  severity failure;
	assert RAM(29689) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(29689))))  severity failure;
	assert RAM(29690) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(29690))))  severity failure;
	assert RAM(29691) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(29691))))  severity failure;
	assert RAM(29692) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29692))))  severity failure;
	assert RAM(29693) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(29693))))  severity failure;
	assert RAM(29694) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(29694))))  severity failure;
	assert RAM(29695) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(29695))))  severity failure;
	assert RAM(29696) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(29696))))  severity failure;
	assert RAM(29697) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29697))))  severity failure;
	assert RAM(29698) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29698))))  severity failure;
	assert RAM(29699) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29699))))  severity failure;
	assert RAM(29700) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(29700))))  severity failure;
	assert RAM(29701) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29701))))  severity failure;
	assert RAM(29702) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29702))))  severity failure;
	assert RAM(29703) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(29703))))  severity failure;
	assert RAM(29704) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(29704))))  severity failure;
	assert RAM(29705) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29705))))  severity failure;
	assert RAM(29706) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(29706))))  severity failure;
	assert RAM(29707) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(29707))))  severity failure;
	assert RAM(29708) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(29708))))  severity failure;
	assert RAM(29709) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(29709))))  severity failure;
	assert RAM(29710) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(29710))))  severity failure;
	assert RAM(29711) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29711))))  severity failure;
	assert RAM(29712) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(29712))))  severity failure;
	assert RAM(29713) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(29713))))  severity failure;
	assert RAM(29714) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(29714))))  severity failure;
	assert RAM(29715) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(29715))))  severity failure;
	assert RAM(29716) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(29716))))  severity failure;
	assert RAM(29717) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(29717))))  severity failure;
	assert RAM(29718) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(29718))))  severity failure;
	assert RAM(29719) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29719))))  severity failure;
	assert RAM(29720) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(29720))))  severity failure;
	assert RAM(29721) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(29721))))  severity failure;
	assert RAM(29722) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(29722))))  severity failure;
	assert RAM(29723) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(29723))))  severity failure;
	assert RAM(29724) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(29724))))  severity failure;
	assert RAM(29725) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(29725))))  severity failure;
	assert RAM(29726) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(29726))))  severity failure;
	assert RAM(29727) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29727))))  severity failure;
	assert RAM(29728) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29728))))  severity failure;
	assert RAM(29729) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(29729))))  severity failure;
	assert RAM(29730) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(29730))))  severity failure;
	assert RAM(29731) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29731))))  severity failure;
	assert RAM(29732) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(29732))))  severity failure;
	assert RAM(29733) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(29733))))  severity failure;
	assert RAM(29734) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29734))))  severity failure;
	assert RAM(29735) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(29735))))  severity failure;
	assert RAM(29736) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29736))))  severity failure;
	assert RAM(29737) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29737))))  severity failure;
	assert RAM(29738) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(29738))))  severity failure;
	assert RAM(29739) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(29739))))  severity failure;
	assert RAM(29740) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29740))))  severity failure;
	assert RAM(29741) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(29741))))  severity failure;
	assert RAM(29742) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(29742))))  severity failure;
	assert RAM(29743) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(29743))))  severity failure;
	assert RAM(29744) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(29744))))  severity failure;
	assert RAM(29745) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(29745))))  severity failure;
	assert RAM(29746) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(29746))))  severity failure;
	assert RAM(29747) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(29747))))  severity failure;
	assert RAM(29748) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(29748))))  severity failure;
	assert RAM(29749) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(29749))))  severity failure;
	assert RAM(29750) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(29750))))  severity failure;
	assert RAM(29751) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(29751))))  severity failure;
	assert RAM(29752) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(29752))))  severity failure;
	assert RAM(29753) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(29753))))  severity failure;
	assert RAM(29754) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(29754))))  severity failure;
	assert RAM(29755) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29755))))  severity failure;
	assert RAM(29756) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(29756))))  severity failure;
	assert RAM(29757) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(29757))))  severity failure;
	assert RAM(29758) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(29758))))  severity failure;
	assert RAM(29759) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(29759))))  severity failure;
	assert RAM(29760) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(29760))))  severity failure;
	assert RAM(29761) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(29761))))  severity failure;
	assert RAM(29762) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(29762))))  severity failure;
	assert RAM(29763) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29763))))  severity failure;
	assert RAM(29764) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(29764))))  severity failure;
	assert RAM(29765) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(29765))))  severity failure;
	assert RAM(29766) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(29766))))  severity failure;
	assert RAM(29767) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(29767))))  severity failure;
	assert RAM(29768) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(29768))))  severity failure;
	assert RAM(29769) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(29769))))  severity failure;
	assert RAM(29770) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(29770))))  severity failure;
	assert RAM(29771) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(29771))))  severity failure;
	assert RAM(29772) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(29772))))  severity failure;
	assert RAM(29773) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(29773))))  severity failure;
	assert RAM(29774) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(29774))))  severity failure;
	assert RAM(29775) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29775))))  severity failure;
	assert RAM(29776) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(29776))))  severity failure;
	assert RAM(29777) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(29777))))  severity failure;
	assert RAM(29778) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(29778))))  severity failure;
	assert RAM(29779) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29779))))  severity failure;
	assert RAM(29780) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29780))))  severity failure;
	assert RAM(29781) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(29781))))  severity failure;
	assert RAM(29782) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(29782))))  severity failure;
	assert RAM(29783) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(29783))))  severity failure;
	assert RAM(29784) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(29784))))  severity failure;
	assert RAM(29785) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(29785))))  severity failure;
	assert RAM(29786) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(29786))))  severity failure;
	assert RAM(29787) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(29787))))  severity failure;
	assert RAM(29788) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(29788))))  severity failure;
	assert RAM(29789) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29789))))  severity failure;
	assert RAM(29790) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29790))))  severity failure;
	assert RAM(29791) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(29791))))  severity failure;
	assert RAM(29792) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29792))))  severity failure;
	assert RAM(29793) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(29793))))  severity failure;
	assert RAM(29794) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(29794))))  severity failure;
	assert RAM(29795) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(29795))))  severity failure;
	assert RAM(29796) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(29796))))  severity failure;
	assert RAM(29797) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29797))))  severity failure;
	assert RAM(29798) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(29798))))  severity failure;
	assert RAM(29799) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(29799))))  severity failure;
	assert RAM(29800) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(29800))))  severity failure;
	assert RAM(29801) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(29801))))  severity failure;
	assert RAM(29802) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29802))))  severity failure;
	assert RAM(29803) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(29803))))  severity failure;
	assert RAM(29804) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(29804))))  severity failure;
	assert RAM(29805) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(29805))))  severity failure;
	assert RAM(29806) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(29806))))  severity failure;
	assert RAM(29807) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29807))))  severity failure;
	assert RAM(29808) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(29808))))  severity failure;
	assert RAM(29809) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29809))))  severity failure;
	assert RAM(29810) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29810))))  severity failure;
	assert RAM(29811) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(29811))))  severity failure;
	assert RAM(29812) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29812))))  severity failure;
	assert RAM(29813) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(29813))))  severity failure;
	assert RAM(29814) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29814))))  severity failure;
	assert RAM(29815) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(29815))))  severity failure;
	assert RAM(29816) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(29816))))  severity failure;
	assert RAM(29817) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(29817))))  severity failure;
	assert RAM(29818) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(29818))))  severity failure;
	assert RAM(29819) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(29819))))  severity failure;
	assert RAM(29820) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(29820))))  severity failure;
	assert RAM(29821) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(29821))))  severity failure;
	assert RAM(29822) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(29822))))  severity failure;
	assert RAM(29823) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(29823))))  severity failure;
	assert RAM(29824) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(29824))))  severity failure;
	assert RAM(29825) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(29825))))  severity failure;
	assert RAM(29826) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(29826))))  severity failure;
	assert RAM(29827) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(29827))))  severity failure;
	assert RAM(29828) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(29828))))  severity failure;
	assert RAM(29829) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(29829))))  severity failure;
	assert RAM(29830) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(29830))))  severity failure;
	assert RAM(29831) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(29831))))  severity failure;
	assert RAM(29832) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(29832))))  severity failure;
	assert RAM(29833) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(29833))))  severity failure;
	assert RAM(29834) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(29834))))  severity failure;
	assert RAM(29835) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29835))))  severity failure;
	assert RAM(29836) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(29836))))  severity failure;
	assert RAM(29837) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29837))))  severity failure;
	assert RAM(29838) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(29838))))  severity failure;
	assert RAM(29839) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(29839))))  severity failure;
	assert RAM(29840) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(29840))))  severity failure;
	assert RAM(29841) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(29841))))  severity failure;
	assert RAM(29842) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29842))))  severity failure;
	assert RAM(29843) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29843))))  severity failure;
	assert RAM(29844) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(29844))))  severity failure;
	assert RAM(29845) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(29845))))  severity failure;
	assert RAM(29846) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(29846))))  severity failure;
	assert RAM(29847) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(29847))))  severity failure;
	assert RAM(29848) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(29848))))  severity failure;
	assert RAM(29849) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(29849))))  severity failure;
	assert RAM(29850) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29850))))  severity failure;
	assert RAM(29851) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(29851))))  severity failure;
	assert RAM(29852) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(29852))))  severity failure;
	assert RAM(29853) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(29853))))  severity failure;
	assert RAM(29854) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29854))))  severity failure;
	assert RAM(29855) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(29855))))  severity failure;
	assert RAM(29856) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(29856))))  severity failure;
	assert RAM(29857) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(29857))))  severity failure;
	assert RAM(29858) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(29858))))  severity failure;
	assert RAM(29859) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(29859))))  severity failure;
	assert RAM(29860) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(29860))))  severity failure;
	assert RAM(29861) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(29861))))  severity failure;
	assert RAM(29862) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(29862))))  severity failure;
	assert RAM(29863) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(29863))))  severity failure;
	assert RAM(29864) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29864))))  severity failure;
	assert RAM(29865) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(29865))))  severity failure;
	assert RAM(29866) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(29866))))  severity failure;
	assert RAM(29867) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(29867))))  severity failure;
	assert RAM(29868) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(29868))))  severity failure;
	assert RAM(29869) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29869))))  severity failure;
	assert RAM(29870) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(29870))))  severity failure;
	assert RAM(29871) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(29871))))  severity failure;
	assert RAM(29872) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(29872))))  severity failure;
	assert RAM(29873) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(29873))))  severity failure;
	assert RAM(29874) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29874))))  severity failure;
	assert RAM(29875) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(29875))))  severity failure;
	assert RAM(29876) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29876))))  severity failure;
	assert RAM(29877) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(29877))))  severity failure;
	assert RAM(29878) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29878))))  severity failure;
	assert RAM(29879) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(29879))))  severity failure;
	assert RAM(29880) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(29880))))  severity failure;
	assert RAM(29881) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29881))))  severity failure;
	assert RAM(29882) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(29882))))  severity failure;
	assert RAM(29883) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29883))))  severity failure;
	assert RAM(29884) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29884))))  severity failure;
	assert RAM(29885) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(29885))))  severity failure;
	assert RAM(29886) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(29886))))  severity failure;
	assert RAM(29887) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(29887))))  severity failure;
	assert RAM(29888) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(29888))))  severity failure;
	assert RAM(29889) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(29889))))  severity failure;
	assert RAM(29890) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(29890))))  severity failure;
	assert RAM(29891) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(29891))))  severity failure;
	assert RAM(29892) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29892))))  severity failure;
	assert RAM(29893) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(29893))))  severity failure;
	assert RAM(29894) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(29894))))  severity failure;
	assert RAM(29895) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29895))))  severity failure;
	assert RAM(29896) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(29896))))  severity failure;
	assert RAM(29897) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(29897))))  severity failure;
	assert RAM(29898) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(29898))))  severity failure;
	assert RAM(29899) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(29899))))  severity failure;
	assert RAM(29900) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(29900))))  severity failure;
	assert RAM(29901) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(29901))))  severity failure;
	assert RAM(29902) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(29902))))  severity failure;
	assert RAM(29903) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(29903))))  severity failure;
	assert RAM(29904) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29904))))  severity failure;
	assert RAM(29905) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(29905))))  severity failure;
	assert RAM(29906) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(29906))))  severity failure;
	assert RAM(29907) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29907))))  severity failure;
	assert RAM(29908) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(29908))))  severity failure;
	assert RAM(29909) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(29909))))  severity failure;
	assert RAM(29910) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(29910))))  severity failure;
	assert RAM(29911) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(29911))))  severity failure;
	assert RAM(29912) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(29912))))  severity failure;
	assert RAM(29913) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(29913))))  severity failure;
	assert RAM(29914) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(29914))))  severity failure;
	assert RAM(29915) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(29915))))  severity failure;
	assert RAM(29916) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(29916))))  severity failure;
	assert RAM(29917) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(29917))))  severity failure;
	assert RAM(29918) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(29918))))  severity failure;
	assert RAM(29919) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(29919))))  severity failure;
	assert RAM(29920) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(29920))))  severity failure;
	assert RAM(29921) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(29921))))  severity failure;
	assert RAM(29922) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(29922))))  severity failure;
	assert RAM(29923) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(29923))))  severity failure;
	assert RAM(29924) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(29924))))  severity failure;
	assert RAM(29925) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29925))))  severity failure;
	assert RAM(29926) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(29926))))  severity failure;
	assert RAM(29927) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29927))))  severity failure;
	assert RAM(29928) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29928))))  severity failure;
	assert RAM(29929) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(29929))))  severity failure;
	assert RAM(29930) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(29930))))  severity failure;
	assert RAM(29931) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(29931))))  severity failure;
	assert RAM(29932) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(29932))))  severity failure;
	assert RAM(29933) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(29933))))  severity failure;
	assert RAM(29934) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(29934))))  severity failure;
	assert RAM(29935) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(29935))))  severity failure;
	assert RAM(29936) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(29936))))  severity failure;
	assert RAM(29937) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29937))))  severity failure;
	assert RAM(29938) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(29938))))  severity failure;
	assert RAM(29939) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(29939))))  severity failure;
	assert RAM(29940) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(29940))))  severity failure;
	assert RAM(29941) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(29941))))  severity failure;
	assert RAM(29942) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(29942))))  severity failure;
	assert RAM(29943) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29943))))  severity failure;
	assert RAM(29944) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(29944))))  severity failure;
	assert RAM(29945) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(29945))))  severity failure;
	assert RAM(29946) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(29946))))  severity failure;
	assert RAM(29947) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(29947))))  severity failure;
	assert RAM(29948) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(29948))))  severity failure;
	assert RAM(29949) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(29949))))  severity failure;
	assert RAM(29950) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(29950))))  severity failure;
	assert RAM(29951) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(29951))))  severity failure;
	assert RAM(29952) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(29952))))  severity failure;
	assert RAM(29953) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(29953))))  severity failure;
	assert RAM(29954) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(29954))))  severity failure;
	assert RAM(29955) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(29955))))  severity failure;
	assert RAM(29956) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(29956))))  severity failure;
	assert RAM(29957) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(29957))))  severity failure;
	assert RAM(29958) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(29958))))  severity failure;
	assert RAM(29959) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(29959))))  severity failure;
	assert RAM(29960) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(29960))))  severity failure;
	assert RAM(29961) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(29961))))  severity failure;
	assert RAM(29962) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(29962))))  severity failure;
	assert RAM(29963) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(29963))))  severity failure;
	assert RAM(29964) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(29964))))  severity failure;
	assert RAM(29965) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(29965))))  severity failure;
	assert RAM(29966) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(29966))))  severity failure;
	assert RAM(29967) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(29967))))  severity failure;
	assert RAM(29968) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(29968))))  severity failure;
	assert RAM(29969) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(29969))))  severity failure;
	assert RAM(29970) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(29970))))  severity failure;
	assert RAM(29971) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(29971))))  severity failure;
	assert RAM(29972) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(29972))))  severity failure;
	assert RAM(29973) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(29973))))  severity failure;
	assert RAM(29974) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(29974))))  severity failure;
	assert RAM(29975) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(29975))))  severity failure;
	assert RAM(29976) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(29976))))  severity failure;
	assert RAM(29977) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(29977))))  severity failure;
	assert RAM(29978) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(29978))))  severity failure;
	assert RAM(29979) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(29979))))  severity failure;
	assert RAM(29980) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(29980))))  severity failure;
	assert RAM(29981) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(29981))))  severity failure;
	assert RAM(29982) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(29982))))  severity failure;
	assert RAM(29983) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(29983))))  severity failure;
	assert RAM(29984) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(29984))))  severity failure;
	assert RAM(29985) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(29985))))  severity failure;
	assert RAM(29986) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(29986))))  severity failure;
	assert RAM(29987) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29987))))  severity failure;
	assert RAM(29988) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(29988))))  severity failure;
	assert RAM(29989) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(29989))))  severity failure;
	assert RAM(29990) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(29990))))  severity failure;
	assert RAM(29991) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(29991))))  severity failure;
	assert RAM(29992) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(29992))))  severity failure;
	assert RAM(29993) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(29993))))  severity failure;
	assert RAM(29994) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(29994))))  severity failure;
	assert RAM(29995) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(29995))))  severity failure;
	assert RAM(29996) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(29996))))  severity failure;
	assert RAM(29997) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29997))))  severity failure;
	assert RAM(29998) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(29998))))  severity failure;
	assert RAM(29999) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(29999))))  severity failure;
	assert RAM(30000) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30000))))  severity failure;
	assert RAM(30001) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(30001))))  severity failure;
	assert RAM(30002) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(30002))))  severity failure;
	assert RAM(30003) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(30003))))  severity failure;
	assert RAM(30004) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30004))))  severity failure;
	assert RAM(30005) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30005))))  severity failure;
	assert RAM(30006) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(30006))))  severity failure;
	assert RAM(30007) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(30007))))  severity failure;
	assert RAM(30008) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(30008))))  severity failure;
	assert RAM(30009) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30009))))  severity failure;
	assert RAM(30010) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30010))))  severity failure;
	assert RAM(30011) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(30011))))  severity failure;
	assert RAM(30012) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(30012))))  severity failure;
	assert RAM(30013) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30013))))  severity failure;
	assert RAM(30014) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(30014))))  severity failure;
	assert RAM(30015) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30015))))  severity failure;
	assert RAM(30016) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(30016))))  severity failure;
	assert RAM(30017) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30017))))  severity failure;
	assert RAM(30018) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30018))))  severity failure;
	assert RAM(30019) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30019))))  severity failure;
	assert RAM(30020) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30020))))  severity failure;
	assert RAM(30021) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(30021))))  severity failure;
	assert RAM(30022) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(30022))))  severity failure;
	assert RAM(30023) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(30023))))  severity failure;
	assert RAM(30024) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(30024))))  severity failure;
	assert RAM(30025) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30025))))  severity failure;
	assert RAM(30026) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(30026))))  severity failure;
	assert RAM(30027) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(30027))))  severity failure;
	assert RAM(30028) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30028))))  severity failure;
	assert RAM(30029) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(30029))))  severity failure;
	assert RAM(30030) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(30030))))  severity failure;
	assert RAM(30031) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(30031))))  severity failure;
	assert RAM(30032) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30032))))  severity failure;
	assert RAM(30033) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(30033))))  severity failure;
	assert RAM(30034) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(30034))))  severity failure;
	assert RAM(30035) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(30035))))  severity failure;
	assert RAM(30036) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(30036))))  severity failure;
	assert RAM(30037) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30037))))  severity failure;
	assert RAM(30038) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(30038))))  severity failure;
	assert RAM(30039) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(30039))))  severity failure;
	assert RAM(30040) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30040))))  severity failure;
	assert RAM(30041) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30041))))  severity failure;
	assert RAM(30042) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(30042))))  severity failure;
	assert RAM(30043) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(30043))))  severity failure;
	assert RAM(30044) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(30044))))  severity failure;
	assert RAM(30045) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30045))))  severity failure;
	assert RAM(30046) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(30046))))  severity failure;
	assert RAM(30047) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30047))))  severity failure;
	assert RAM(30048) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(30048))))  severity failure;
	assert RAM(30049) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(30049))))  severity failure;
	assert RAM(30050) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30050))))  severity failure;
	assert RAM(30051) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(30051))))  severity failure;
	assert RAM(30052) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(30052))))  severity failure;
	assert RAM(30053) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(30053))))  severity failure;
	assert RAM(30054) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(30054))))  severity failure;
	assert RAM(30055) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(30055))))  severity failure;
	assert RAM(30056) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30056))))  severity failure;
	assert RAM(30057) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30057))))  severity failure;
	assert RAM(30058) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(30058))))  severity failure;
	assert RAM(30059) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30059))))  severity failure;
	assert RAM(30060) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(30060))))  severity failure;
	assert RAM(30061) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30061))))  severity failure;
	assert RAM(30062) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(30062))))  severity failure;
	assert RAM(30063) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(30063))))  severity failure;
	assert RAM(30064) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(30064))))  severity failure;
	assert RAM(30065) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30065))))  severity failure;
	assert RAM(30066) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(30066))))  severity failure;
	assert RAM(30067) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30067))))  severity failure;
	assert RAM(30068) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(30068))))  severity failure;
	assert RAM(30069) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(30069))))  severity failure;
	assert RAM(30070) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30070))))  severity failure;
	assert RAM(30071) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(30071))))  severity failure;
	assert RAM(30072) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(30072))))  severity failure;
	assert RAM(30073) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30073))))  severity failure;
	assert RAM(30074) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30074))))  severity failure;
	assert RAM(30075) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30075))))  severity failure;
	assert RAM(30076) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30076))))  severity failure;
	assert RAM(30077) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(30077))))  severity failure;
	assert RAM(30078) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(30078))))  severity failure;
	assert RAM(30079) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(30079))))  severity failure;
	assert RAM(30080) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(30080))))  severity failure;
	assert RAM(30081) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30081))))  severity failure;
	assert RAM(30082) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30082))))  severity failure;
	assert RAM(30083) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(30083))))  severity failure;
	assert RAM(30084) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30084))))  severity failure;
	assert RAM(30085) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(30085))))  severity failure;
	assert RAM(30086) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(30086))))  severity failure;
	assert RAM(30087) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(30087))))  severity failure;
	assert RAM(30088) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30088))))  severity failure;
	assert RAM(30089) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(30089))))  severity failure;
	assert RAM(30090) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30090))))  severity failure;
	assert RAM(30091) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(30091))))  severity failure;
	assert RAM(30092) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30092))))  severity failure;
	assert RAM(30093) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30093))))  severity failure;
	assert RAM(30094) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(30094))))  severity failure;
	assert RAM(30095) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(30095))))  severity failure;
	assert RAM(30096) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(30096))))  severity failure;
	assert RAM(30097) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30097))))  severity failure;
	assert RAM(30098) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30098))))  severity failure;
	assert RAM(30099) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(30099))))  severity failure;
	assert RAM(30100) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30100))))  severity failure;
	assert RAM(30101) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(30101))))  severity failure;
	assert RAM(30102) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(30102))))  severity failure;
	assert RAM(30103) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30103))))  severity failure;
	assert RAM(30104) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(30104))))  severity failure;
	assert RAM(30105) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(30105))))  severity failure;
	assert RAM(30106) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30106))))  severity failure;
	assert RAM(30107) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(30107))))  severity failure;
	assert RAM(30108) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(30108))))  severity failure;
	assert RAM(30109) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30109))))  severity failure;
	assert RAM(30110) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(30110))))  severity failure;
	assert RAM(30111) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30111))))  severity failure;
	assert RAM(30112) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30112))))  severity failure;
	assert RAM(30113) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(30113))))  severity failure;
	assert RAM(30114) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(30114))))  severity failure;
	assert RAM(30115) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(30115))))  severity failure;
	assert RAM(30116) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(30116))))  severity failure;
	assert RAM(30117) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30117))))  severity failure;
	assert RAM(30118) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(30118))))  severity failure;
	assert RAM(30119) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(30119))))  severity failure;
	assert RAM(30120) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30120))))  severity failure;
	assert RAM(30121) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30121))))  severity failure;
	assert RAM(30122) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30122))))  severity failure;
	assert RAM(30123) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(30123))))  severity failure;
	assert RAM(30124) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(30124))))  severity failure;
	assert RAM(30125) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30125))))  severity failure;
	assert RAM(30126) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(30126))))  severity failure;
	assert RAM(30127) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(30127))))  severity failure;
	assert RAM(30128) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(30128))))  severity failure;
	assert RAM(30129) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(30129))))  severity failure;
	assert RAM(30130) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(30130))))  severity failure;
	assert RAM(30131) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(30131))))  severity failure;
	assert RAM(30132) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(30132))))  severity failure;
	assert RAM(30133) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(30133))))  severity failure;
	assert RAM(30134) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30134))))  severity failure;
	assert RAM(30135) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30135))))  severity failure;
	assert RAM(30136) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30136))))  severity failure;
	assert RAM(30137) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(30137))))  severity failure;
	assert RAM(30138) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30138))))  severity failure;
	assert RAM(30139) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(30139))))  severity failure;
	assert RAM(30140) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(30140))))  severity failure;
	assert RAM(30141) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(30141))))  severity failure;
	assert RAM(30142) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30142))))  severity failure;
	assert RAM(30143) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(30143))))  severity failure;
	assert RAM(30144) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(30144))))  severity failure;
	assert RAM(30145) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30145))))  severity failure;
	assert RAM(30146) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30146))))  severity failure;
	assert RAM(30147) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30147))))  severity failure;
	assert RAM(30148) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30148))))  severity failure;
	assert RAM(30149) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(30149))))  severity failure;
	assert RAM(30150) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(30150))))  severity failure;
	assert RAM(30151) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(30151))))  severity failure;
	assert RAM(30152) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(30152))))  severity failure;
	assert RAM(30153) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30153))))  severity failure;
	assert RAM(30154) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(30154))))  severity failure;
	assert RAM(30155) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30155))))  severity failure;
	assert RAM(30156) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(30156))))  severity failure;
	assert RAM(30157) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(30157))))  severity failure;
	assert RAM(30158) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(30158))))  severity failure;
	assert RAM(30159) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(30159))))  severity failure;
	assert RAM(30160) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(30160))))  severity failure;
	assert RAM(30161) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(30161))))  severity failure;
	assert RAM(30162) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30162))))  severity failure;
	assert RAM(30163) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30163))))  severity failure;
	assert RAM(30164) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(30164))))  severity failure;
	assert RAM(30165) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30165))))  severity failure;
	assert RAM(30166) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(30166))))  severity failure;
	assert RAM(30167) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30167))))  severity failure;
	assert RAM(30168) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(30168))))  severity failure;
	assert RAM(30169) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(30169))))  severity failure;
	assert RAM(30170) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30170))))  severity failure;
	assert RAM(30171) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(30171))))  severity failure;
	assert RAM(30172) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30172))))  severity failure;
	assert RAM(30173) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(30173))))  severity failure;
	assert RAM(30174) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(30174))))  severity failure;
	assert RAM(30175) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(30175))))  severity failure;
	assert RAM(30176) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30176))))  severity failure;
	assert RAM(30177) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(30177))))  severity failure;
	assert RAM(30178) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30178))))  severity failure;
	assert RAM(30179) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(30179))))  severity failure;
	assert RAM(30180) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(30180))))  severity failure;
	assert RAM(30181) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(30181))))  severity failure;
	assert RAM(30182) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(30182))))  severity failure;
	assert RAM(30183) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30183))))  severity failure;
	assert RAM(30184) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(30184))))  severity failure;
	assert RAM(30185) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(30185))))  severity failure;
	assert RAM(30186) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30186))))  severity failure;
	assert RAM(30187) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(30187))))  severity failure;
	assert RAM(30188) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30188))))  severity failure;
	assert RAM(30189) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(30189))))  severity failure;
	assert RAM(30190) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(30190))))  severity failure;
	assert RAM(30191) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30191))))  severity failure;
	assert RAM(30192) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(30192))))  severity failure;
	assert RAM(30193) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30193))))  severity failure;
	assert RAM(30194) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30194))))  severity failure;
	assert RAM(30195) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(30195))))  severity failure;
	assert RAM(30196) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(30196))))  severity failure;
	assert RAM(30197) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30197))))  severity failure;
	assert RAM(30198) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30198))))  severity failure;
	assert RAM(30199) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30199))))  severity failure;
	assert RAM(30200) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(30200))))  severity failure;
	assert RAM(30201) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(30201))))  severity failure;
	assert RAM(30202) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30202))))  severity failure;
	assert RAM(30203) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(30203))))  severity failure;
	assert RAM(30204) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(30204))))  severity failure;
	assert RAM(30205) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(30205))))  severity failure;
	assert RAM(30206) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(30206))))  severity failure;
	assert RAM(30207) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30207))))  severity failure;
	assert RAM(30208) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30208))))  severity failure;
	assert RAM(30209) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(30209))))  severity failure;
	assert RAM(30210) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30210))))  severity failure;
	assert RAM(30211) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(30211))))  severity failure;
	assert RAM(30212) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(30212))))  severity failure;
	assert RAM(30213) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30213))))  severity failure;
	assert RAM(30214) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(30214))))  severity failure;
	assert RAM(30215) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(30215))))  severity failure;
	assert RAM(30216) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(30216))))  severity failure;
	assert RAM(30217) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(30217))))  severity failure;
	assert RAM(30218) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(30218))))  severity failure;
	assert RAM(30219) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30219))))  severity failure;
	assert RAM(30220) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(30220))))  severity failure;
	assert RAM(30221) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(30221))))  severity failure;
	assert RAM(30222) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(30222))))  severity failure;
	assert RAM(30223) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30223))))  severity failure;
	assert RAM(30224) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(30224))))  severity failure;
	assert RAM(30225) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(30225))))  severity failure;
	assert RAM(30226) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(30226))))  severity failure;
	assert RAM(30227) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(30227))))  severity failure;
	assert RAM(30228) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(30228))))  severity failure;
	assert RAM(30229) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30229))))  severity failure;
	assert RAM(30230) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(30230))))  severity failure;
	assert RAM(30231) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(30231))))  severity failure;
	assert RAM(30232) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(30232))))  severity failure;
	assert RAM(30233) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30233))))  severity failure;
	assert RAM(30234) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(30234))))  severity failure;
	assert RAM(30235) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(30235))))  severity failure;
	assert RAM(30236) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(30236))))  severity failure;
	assert RAM(30237) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(30237))))  severity failure;
	assert RAM(30238) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30238))))  severity failure;
	assert RAM(30239) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30239))))  severity failure;
	assert RAM(30240) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30240))))  severity failure;
	assert RAM(30241) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30241))))  severity failure;
	assert RAM(30242) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30242))))  severity failure;
	assert RAM(30243) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30243))))  severity failure;
	assert RAM(30244) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(30244))))  severity failure;
	assert RAM(30245) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(30245))))  severity failure;
	assert RAM(30246) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30246))))  severity failure;
	assert RAM(30247) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(30247))))  severity failure;
	assert RAM(30248) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(30248))))  severity failure;
	assert RAM(30249) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(30249))))  severity failure;
	assert RAM(30250) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(30250))))  severity failure;
	assert RAM(30251) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30251))))  severity failure;
	assert RAM(30252) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30252))))  severity failure;
	assert RAM(30253) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(30253))))  severity failure;
	assert RAM(30254) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(30254))))  severity failure;
	assert RAM(30255) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(30255))))  severity failure;
	assert RAM(30256) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(30256))))  severity failure;
	assert RAM(30257) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30257))))  severity failure;
	assert RAM(30258) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(30258))))  severity failure;
	assert RAM(30259) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30259))))  severity failure;
	assert RAM(30260) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30260))))  severity failure;
	assert RAM(30261) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30261))))  severity failure;
	assert RAM(30262) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30262))))  severity failure;
	assert RAM(30263) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30263))))  severity failure;
	assert RAM(30264) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(30264))))  severity failure;
	assert RAM(30265) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30265))))  severity failure;
	assert RAM(30266) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30266))))  severity failure;
	assert RAM(30267) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(30267))))  severity failure;
	assert RAM(30268) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(30268))))  severity failure;
	assert RAM(30269) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30269))))  severity failure;
	assert RAM(30270) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(30270))))  severity failure;
	assert RAM(30271) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30271))))  severity failure;
	assert RAM(30272) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30272))))  severity failure;
	assert RAM(30273) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(30273))))  severity failure;
	assert RAM(30274) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(30274))))  severity failure;
	assert RAM(30275) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(30275))))  severity failure;
	assert RAM(30276) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(30276))))  severity failure;
	assert RAM(30277) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(30277))))  severity failure;
	assert RAM(30278) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(30278))))  severity failure;
	assert RAM(30279) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30279))))  severity failure;
	assert RAM(30280) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(30280))))  severity failure;
	assert RAM(30281) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(30281))))  severity failure;
	assert RAM(30282) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30282))))  severity failure;
	assert RAM(30283) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(30283))))  severity failure;
	assert RAM(30284) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(30284))))  severity failure;
	assert RAM(30285) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(30285))))  severity failure;
	assert RAM(30286) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(30286))))  severity failure;
	assert RAM(30287) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30287))))  severity failure;
	assert RAM(30288) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30288))))  severity failure;
	assert RAM(30289) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30289))))  severity failure;
	assert RAM(30290) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(30290))))  severity failure;
	assert RAM(30291) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30291))))  severity failure;
	assert RAM(30292) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30292))))  severity failure;
	assert RAM(30293) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(30293))))  severity failure;
	assert RAM(30294) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(30294))))  severity failure;
	assert RAM(30295) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(30295))))  severity failure;
	assert RAM(30296) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(30296))))  severity failure;
	assert RAM(30297) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(30297))))  severity failure;
	assert RAM(30298) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(30298))))  severity failure;
	assert RAM(30299) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30299))))  severity failure;
	assert RAM(30300) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(30300))))  severity failure;
	assert RAM(30301) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30301))))  severity failure;
	assert RAM(30302) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30302))))  severity failure;
	assert RAM(30303) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30303))))  severity failure;
	assert RAM(30304) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(30304))))  severity failure;
	assert RAM(30305) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(30305))))  severity failure;
	assert RAM(30306) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30306))))  severity failure;
	assert RAM(30307) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(30307))))  severity failure;
	assert RAM(30308) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(30308))))  severity failure;
	assert RAM(30309) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(30309))))  severity failure;
	assert RAM(30310) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30310))))  severity failure;
	assert RAM(30311) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30311))))  severity failure;
	assert RAM(30312) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30312))))  severity failure;
	assert RAM(30313) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30313))))  severity failure;
	assert RAM(30314) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(30314))))  severity failure;
	assert RAM(30315) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(30315))))  severity failure;
	assert RAM(30316) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(30316))))  severity failure;
	assert RAM(30317) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(30317))))  severity failure;
	assert RAM(30318) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30318))))  severity failure;
	assert RAM(30319) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(30319))))  severity failure;
	assert RAM(30320) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(30320))))  severity failure;
	assert RAM(30321) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30321))))  severity failure;
	assert RAM(30322) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(30322))))  severity failure;
	assert RAM(30323) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(30323))))  severity failure;
	assert RAM(30324) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(30324))))  severity failure;
	assert RAM(30325) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(30325))))  severity failure;
	assert RAM(30326) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(30326))))  severity failure;
	assert RAM(30327) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30327))))  severity failure;
	assert RAM(30328) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(30328))))  severity failure;
	assert RAM(30329) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(30329))))  severity failure;
	assert RAM(30330) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30330))))  severity failure;
	assert RAM(30331) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(30331))))  severity failure;
	assert RAM(30332) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(30332))))  severity failure;
	assert RAM(30333) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(30333))))  severity failure;
	assert RAM(30334) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(30334))))  severity failure;
	assert RAM(30335) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30335))))  severity failure;
	assert RAM(30336) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30336))))  severity failure;
	assert RAM(30337) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(30337))))  severity failure;
	assert RAM(30338) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(30338))))  severity failure;
	assert RAM(30339) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30339))))  severity failure;
	assert RAM(30340) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30340))))  severity failure;
	assert RAM(30341) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(30341))))  severity failure;
	assert RAM(30342) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(30342))))  severity failure;
	assert RAM(30343) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(30343))))  severity failure;
	assert RAM(30344) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(30344))))  severity failure;
	assert RAM(30345) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30345))))  severity failure;
	assert RAM(30346) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(30346))))  severity failure;
	assert RAM(30347) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30347))))  severity failure;
	assert RAM(30348) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(30348))))  severity failure;
	assert RAM(30349) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(30349))))  severity failure;
	assert RAM(30350) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30350))))  severity failure;
	assert RAM(30351) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(30351))))  severity failure;
	assert RAM(30352) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30352))))  severity failure;
	assert RAM(30353) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30353))))  severity failure;
	assert RAM(30354) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(30354))))  severity failure;
	assert RAM(30355) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(30355))))  severity failure;
	assert RAM(30356) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(30356))))  severity failure;
	assert RAM(30357) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30357))))  severity failure;
	assert RAM(30358) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(30358))))  severity failure;
	assert RAM(30359) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30359))))  severity failure;
	assert RAM(30360) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30360))))  severity failure;
	assert RAM(30361) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(30361))))  severity failure;
	assert RAM(30362) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(30362))))  severity failure;
	assert RAM(30363) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(30363))))  severity failure;
	assert RAM(30364) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30364))))  severity failure;
	assert RAM(30365) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30365))))  severity failure;
	assert RAM(30366) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30366))))  severity failure;
	assert RAM(30367) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(30367))))  severity failure;
	assert RAM(30368) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(30368))))  severity failure;
	assert RAM(30369) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30369))))  severity failure;
	assert RAM(30370) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(30370))))  severity failure;
	assert RAM(30371) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(30371))))  severity failure;
	assert RAM(30372) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30372))))  severity failure;
	assert RAM(30373) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30373))))  severity failure;
	assert RAM(30374) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(30374))))  severity failure;
	assert RAM(30375) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30375))))  severity failure;
	assert RAM(30376) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(30376))))  severity failure;
	assert RAM(30377) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30377))))  severity failure;
	assert RAM(30378) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(30378))))  severity failure;
	assert RAM(30379) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(30379))))  severity failure;
	assert RAM(30380) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(30380))))  severity failure;
	assert RAM(30381) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(30381))))  severity failure;
	assert RAM(30382) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(30382))))  severity failure;
	assert RAM(30383) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(30383))))  severity failure;
	assert RAM(30384) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(30384))))  severity failure;
	assert RAM(30385) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(30385))))  severity failure;
	assert RAM(30386) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(30386))))  severity failure;
	assert RAM(30387) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(30387))))  severity failure;
	assert RAM(30388) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(30388))))  severity failure;
	assert RAM(30389) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30389))))  severity failure;
	assert RAM(30390) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(30390))))  severity failure;
	assert RAM(30391) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(30391))))  severity failure;
	assert RAM(30392) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(30392))))  severity failure;
	assert RAM(30393) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(30393))))  severity failure;
	assert RAM(30394) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30394))))  severity failure;
	assert RAM(30395) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(30395))))  severity failure;
	assert RAM(30396) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(30396))))  severity failure;
	assert RAM(30397) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30397))))  severity failure;
	assert RAM(30398) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30398))))  severity failure;
	assert RAM(30399) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30399))))  severity failure;
	assert RAM(30400) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(30400))))  severity failure;
	assert RAM(30401) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30401))))  severity failure;
	assert RAM(30402) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30402))))  severity failure;
	assert RAM(30403) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30403))))  severity failure;
	assert RAM(30404) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30404))))  severity failure;
	assert RAM(30405) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(30405))))  severity failure;
	assert RAM(30406) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30406))))  severity failure;
	assert RAM(30407) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30407))))  severity failure;
	assert RAM(30408) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(30408))))  severity failure;
	assert RAM(30409) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30409))))  severity failure;
	assert RAM(30410) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(30410))))  severity failure;
	assert RAM(30411) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(30411))))  severity failure;
	assert RAM(30412) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(30412))))  severity failure;
	assert RAM(30413) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(30413))))  severity failure;
	assert RAM(30414) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(30414))))  severity failure;
	assert RAM(30415) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30415))))  severity failure;
	assert RAM(30416) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(30416))))  severity failure;
	assert RAM(30417) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(30417))))  severity failure;
	assert RAM(30418) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30418))))  severity failure;
	assert RAM(30419) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(30419))))  severity failure;
	assert RAM(30420) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30420))))  severity failure;
	assert RAM(30421) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(30421))))  severity failure;
	assert RAM(30422) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(30422))))  severity failure;
	assert RAM(30423) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30423))))  severity failure;
	assert RAM(30424) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30424))))  severity failure;
	assert RAM(30425) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(30425))))  severity failure;
	assert RAM(30426) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(30426))))  severity failure;
	assert RAM(30427) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30427))))  severity failure;
	assert RAM(30428) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30428))))  severity failure;
	assert RAM(30429) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30429))))  severity failure;
	assert RAM(30430) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30430))))  severity failure;
	assert RAM(30431) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30431))))  severity failure;
	assert RAM(30432) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(30432))))  severity failure;
	assert RAM(30433) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(30433))))  severity failure;
	assert RAM(30434) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(30434))))  severity failure;
	assert RAM(30435) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(30435))))  severity failure;
	assert RAM(30436) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(30436))))  severity failure;
	assert RAM(30437) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30437))))  severity failure;
	assert RAM(30438) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(30438))))  severity failure;
	assert RAM(30439) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(30439))))  severity failure;
	assert RAM(30440) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30440))))  severity failure;
	assert RAM(30441) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(30441))))  severity failure;
	assert RAM(30442) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(30442))))  severity failure;
	assert RAM(30443) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(30443))))  severity failure;
	assert RAM(30444) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30444))))  severity failure;
	assert RAM(30445) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(30445))))  severity failure;
	assert RAM(30446) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(30446))))  severity failure;
	assert RAM(30447) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(30447))))  severity failure;
	assert RAM(30448) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30448))))  severity failure;
	assert RAM(30449) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(30449))))  severity failure;
	assert RAM(30450) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(30450))))  severity failure;
	assert RAM(30451) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30451))))  severity failure;
	assert RAM(30452) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30452))))  severity failure;
	assert RAM(30453) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(30453))))  severity failure;
	assert RAM(30454) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(30454))))  severity failure;
	assert RAM(30455) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(30455))))  severity failure;
	assert RAM(30456) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30456))))  severity failure;
	assert RAM(30457) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(30457))))  severity failure;
	assert RAM(30458) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(30458))))  severity failure;
	assert RAM(30459) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30459))))  severity failure;
	assert RAM(30460) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(30460))))  severity failure;
	assert RAM(30461) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30461))))  severity failure;
	assert RAM(30462) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(30462))))  severity failure;
	assert RAM(30463) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(30463))))  severity failure;
	assert RAM(30464) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(30464))))  severity failure;
	assert RAM(30465) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(30465))))  severity failure;
	assert RAM(30466) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30466))))  severity failure;
	assert RAM(30467) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(30467))))  severity failure;
	assert RAM(30468) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30468))))  severity failure;
	assert RAM(30469) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(30469))))  severity failure;
	assert RAM(30470) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(30470))))  severity failure;
	assert RAM(30471) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(30471))))  severity failure;
	assert RAM(30472) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(30472))))  severity failure;
	assert RAM(30473) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30473))))  severity failure;
	assert RAM(30474) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30474))))  severity failure;
	assert RAM(30475) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(30475))))  severity failure;
	assert RAM(30476) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(30476))))  severity failure;
	assert RAM(30477) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30477))))  severity failure;
	assert RAM(30478) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(30478))))  severity failure;
	assert RAM(30479) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(30479))))  severity failure;
	assert RAM(30480) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30480))))  severity failure;
	assert RAM(30481) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(30481))))  severity failure;
	assert RAM(30482) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(30482))))  severity failure;
	assert RAM(30483) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(30483))))  severity failure;
	assert RAM(30484) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30484))))  severity failure;
	assert RAM(30485) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(30485))))  severity failure;
	assert RAM(30486) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(30486))))  severity failure;
	assert RAM(30487) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(30487))))  severity failure;
	assert RAM(30488) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(30488))))  severity failure;
	assert RAM(30489) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30489))))  severity failure;
	assert RAM(30490) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(30490))))  severity failure;
	assert RAM(30491) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(30491))))  severity failure;
	assert RAM(30492) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(30492))))  severity failure;
	assert RAM(30493) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30493))))  severity failure;
	assert RAM(30494) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(30494))))  severity failure;
	assert RAM(30495) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(30495))))  severity failure;
	assert RAM(30496) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(30496))))  severity failure;
	assert RAM(30497) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(30497))))  severity failure;
	assert RAM(30498) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(30498))))  severity failure;
	assert RAM(30499) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(30499))))  severity failure;
	assert RAM(30500) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30500))))  severity failure;
	assert RAM(30501) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30501))))  severity failure;
	assert RAM(30502) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30502))))  severity failure;
	assert RAM(30503) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(30503))))  severity failure;
	assert RAM(30504) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30504))))  severity failure;
	assert RAM(30505) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(30505))))  severity failure;
	assert RAM(30506) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30506))))  severity failure;
	assert RAM(30507) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(30507))))  severity failure;
	assert RAM(30508) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30508))))  severity failure;
	assert RAM(30509) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30509))))  severity failure;
	assert RAM(30510) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30510))))  severity failure;
	assert RAM(30511) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30511))))  severity failure;
	assert RAM(30512) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30512))))  severity failure;
	assert RAM(30513) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(30513))))  severity failure;
	assert RAM(30514) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(30514))))  severity failure;
	assert RAM(30515) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(30515))))  severity failure;
	assert RAM(30516) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30516))))  severity failure;
	assert RAM(30517) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(30517))))  severity failure;
	assert RAM(30518) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(30518))))  severity failure;
	assert RAM(30519) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(30519))))  severity failure;
	assert RAM(30520) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(30520))))  severity failure;
	assert RAM(30521) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(30521))))  severity failure;
	assert RAM(30522) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30522))))  severity failure;
	assert RAM(30523) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(30523))))  severity failure;
	assert RAM(30524) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30524))))  severity failure;
	assert RAM(30525) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(30525))))  severity failure;
	assert RAM(30526) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(30526))))  severity failure;
	assert RAM(30527) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(30527))))  severity failure;
	assert RAM(30528) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(30528))))  severity failure;
	assert RAM(30529) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(30529))))  severity failure;
	assert RAM(30530) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30530))))  severity failure;
	assert RAM(30531) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(30531))))  severity failure;
	assert RAM(30532) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30532))))  severity failure;
	assert RAM(30533) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30533))))  severity failure;
	assert RAM(30534) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(30534))))  severity failure;
	assert RAM(30535) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30535))))  severity failure;
	assert RAM(30536) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30536))))  severity failure;
	assert RAM(30537) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(30537))))  severity failure;
	assert RAM(30538) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30538))))  severity failure;
	assert RAM(30539) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(30539))))  severity failure;
	assert RAM(30540) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30540))))  severity failure;
	assert RAM(30541) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(30541))))  severity failure;
	assert RAM(30542) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(30542))))  severity failure;
	assert RAM(30543) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(30543))))  severity failure;
	assert RAM(30544) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(30544))))  severity failure;
	assert RAM(30545) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30545))))  severity failure;
	assert RAM(30546) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30546))))  severity failure;
	assert RAM(30547) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(30547))))  severity failure;
	assert RAM(30548) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30548))))  severity failure;
	assert RAM(30549) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(30549))))  severity failure;
	assert RAM(30550) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30550))))  severity failure;
	assert RAM(30551) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30551))))  severity failure;
	assert RAM(30552) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(30552))))  severity failure;
	assert RAM(30553) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(30553))))  severity failure;
	assert RAM(30554) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(30554))))  severity failure;
	assert RAM(30555) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(30555))))  severity failure;
	assert RAM(30556) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(30556))))  severity failure;
	assert RAM(30557) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30557))))  severity failure;
	assert RAM(30558) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(30558))))  severity failure;
	assert RAM(30559) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30559))))  severity failure;
	assert RAM(30560) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30560))))  severity failure;
	assert RAM(30561) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(30561))))  severity failure;
	assert RAM(30562) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30562))))  severity failure;
	assert RAM(30563) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30563))))  severity failure;
	assert RAM(30564) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(30564))))  severity failure;
	assert RAM(30565) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(30565))))  severity failure;
	assert RAM(30566) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30566))))  severity failure;
	assert RAM(30567) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(30567))))  severity failure;
	assert RAM(30568) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(30568))))  severity failure;
	assert RAM(30569) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30569))))  severity failure;
	assert RAM(30570) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30570))))  severity failure;
	assert RAM(30571) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(30571))))  severity failure;
	assert RAM(30572) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30572))))  severity failure;
	assert RAM(30573) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30573))))  severity failure;
	assert RAM(30574) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30574))))  severity failure;
	assert RAM(30575) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(30575))))  severity failure;
	assert RAM(30576) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(30576))))  severity failure;
	assert RAM(30577) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30577))))  severity failure;
	assert RAM(30578) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(30578))))  severity failure;
	assert RAM(30579) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30579))))  severity failure;
	assert RAM(30580) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(30580))))  severity failure;
	assert RAM(30581) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30581))))  severity failure;
	assert RAM(30582) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(30582))))  severity failure;
	assert RAM(30583) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30583))))  severity failure;
	assert RAM(30584) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(30584))))  severity failure;
	assert RAM(30585) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(30585))))  severity failure;
	assert RAM(30586) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30586))))  severity failure;
	assert RAM(30587) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(30587))))  severity failure;
	assert RAM(30588) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30588))))  severity failure;
	assert RAM(30589) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30589))))  severity failure;
	assert RAM(30590) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(30590))))  severity failure;
	assert RAM(30591) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(30591))))  severity failure;
	assert RAM(30592) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(30592))))  severity failure;
	assert RAM(30593) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30593))))  severity failure;
	assert RAM(30594) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30594))))  severity failure;
	assert RAM(30595) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(30595))))  severity failure;
	assert RAM(30596) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(30596))))  severity failure;
	assert RAM(30597) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(30597))))  severity failure;
	assert RAM(30598) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(30598))))  severity failure;
	assert RAM(30599) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(30599))))  severity failure;
	assert RAM(30600) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(30600))))  severity failure;
	assert RAM(30601) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(30601))))  severity failure;
	assert RAM(30602) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(30602))))  severity failure;
	assert RAM(30603) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30603))))  severity failure;
	assert RAM(30604) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30604))))  severity failure;
	assert RAM(30605) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30605))))  severity failure;
	assert RAM(30606) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(30606))))  severity failure;
	assert RAM(30607) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(30607))))  severity failure;
	assert RAM(30608) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(30608))))  severity failure;
	assert RAM(30609) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30609))))  severity failure;
	assert RAM(30610) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(30610))))  severity failure;
	assert RAM(30611) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30611))))  severity failure;
	assert RAM(30612) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(30612))))  severity failure;
	assert RAM(30613) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30613))))  severity failure;
	assert RAM(30614) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(30614))))  severity failure;
	assert RAM(30615) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30615))))  severity failure;
	assert RAM(30616) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(30616))))  severity failure;
	assert RAM(30617) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(30617))))  severity failure;
	assert RAM(30618) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(30618))))  severity failure;
	assert RAM(30619) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30619))))  severity failure;
	assert RAM(30620) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(30620))))  severity failure;
	assert RAM(30621) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(30621))))  severity failure;
	assert RAM(30622) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(30622))))  severity failure;
	assert RAM(30623) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(30623))))  severity failure;
	assert RAM(30624) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(30624))))  severity failure;
	assert RAM(30625) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(30625))))  severity failure;
	assert RAM(30626) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30626))))  severity failure;
	assert RAM(30627) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30627))))  severity failure;
	assert RAM(30628) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30628))))  severity failure;
	assert RAM(30629) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30629))))  severity failure;
	assert RAM(30630) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(30630))))  severity failure;
	assert RAM(30631) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(30631))))  severity failure;
	assert RAM(30632) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(30632))))  severity failure;
	assert RAM(30633) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(30633))))  severity failure;
	assert RAM(30634) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30634))))  severity failure;
	assert RAM(30635) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(30635))))  severity failure;
	assert RAM(30636) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(30636))))  severity failure;
	assert RAM(30637) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30637))))  severity failure;
	assert RAM(30638) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(30638))))  severity failure;
	assert RAM(30639) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30639))))  severity failure;
	assert RAM(30640) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30640))))  severity failure;
	assert RAM(30641) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(30641))))  severity failure;
	assert RAM(30642) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(30642))))  severity failure;
	assert RAM(30643) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(30643))))  severity failure;
	assert RAM(30644) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30644))))  severity failure;
	assert RAM(30645) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(30645))))  severity failure;
	assert RAM(30646) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30646))))  severity failure;
	assert RAM(30647) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(30647))))  severity failure;
	assert RAM(30648) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30648))))  severity failure;
	assert RAM(30649) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(30649))))  severity failure;
	assert RAM(30650) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(30650))))  severity failure;
	assert RAM(30651) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(30651))))  severity failure;
	assert RAM(30652) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30652))))  severity failure;
	assert RAM(30653) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(30653))))  severity failure;
	assert RAM(30654) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(30654))))  severity failure;
	assert RAM(30655) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(30655))))  severity failure;
	assert RAM(30656) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(30656))))  severity failure;
	assert RAM(30657) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(30657))))  severity failure;
	assert RAM(30658) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(30658))))  severity failure;
	assert RAM(30659) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(30659))))  severity failure;
	assert RAM(30660) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(30660))))  severity failure;
	assert RAM(30661) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30661))))  severity failure;
	assert RAM(30662) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(30662))))  severity failure;
	assert RAM(30663) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(30663))))  severity failure;
	assert RAM(30664) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30664))))  severity failure;
	assert RAM(30665) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(30665))))  severity failure;
	assert RAM(30666) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30666))))  severity failure;
	assert RAM(30667) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(30667))))  severity failure;
	assert RAM(30668) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30668))))  severity failure;
	assert RAM(30669) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(30669))))  severity failure;
	assert RAM(30670) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(30670))))  severity failure;
	assert RAM(30671) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(30671))))  severity failure;
	assert RAM(30672) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(30672))))  severity failure;
	assert RAM(30673) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30673))))  severity failure;
	assert RAM(30674) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(30674))))  severity failure;
	assert RAM(30675) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(30675))))  severity failure;
	assert RAM(30676) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(30676))))  severity failure;
	assert RAM(30677) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(30677))))  severity failure;
	assert RAM(30678) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(30678))))  severity failure;
	assert RAM(30679) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30679))))  severity failure;
	assert RAM(30680) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(30680))))  severity failure;
	assert RAM(30681) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30681))))  severity failure;
	assert RAM(30682) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(30682))))  severity failure;
	assert RAM(30683) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30683))))  severity failure;
	assert RAM(30684) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30684))))  severity failure;
	assert RAM(30685) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(30685))))  severity failure;
	assert RAM(30686) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(30686))))  severity failure;
	assert RAM(30687) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30687))))  severity failure;
	assert RAM(30688) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(30688))))  severity failure;
	assert RAM(30689) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(30689))))  severity failure;
	assert RAM(30690) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(30690))))  severity failure;
	assert RAM(30691) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(30691))))  severity failure;
	assert RAM(30692) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(30692))))  severity failure;
	assert RAM(30693) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(30693))))  severity failure;
	assert RAM(30694) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30694))))  severity failure;
	assert RAM(30695) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(30695))))  severity failure;
	assert RAM(30696) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(30696))))  severity failure;
	assert RAM(30697) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(30697))))  severity failure;
	assert RAM(30698) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(30698))))  severity failure;
	assert RAM(30699) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30699))))  severity failure;
	assert RAM(30700) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(30700))))  severity failure;
	assert RAM(30701) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(30701))))  severity failure;
	assert RAM(30702) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(30702))))  severity failure;
	assert RAM(30703) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(30703))))  severity failure;
	assert RAM(30704) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(30704))))  severity failure;
	assert RAM(30705) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(30705))))  severity failure;
	assert RAM(30706) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(30706))))  severity failure;
	assert RAM(30707) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(30707))))  severity failure;
	assert RAM(30708) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(30708))))  severity failure;
	assert RAM(30709) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(30709))))  severity failure;
	assert RAM(30710) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(30710))))  severity failure;
	assert RAM(30711) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(30711))))  severity failure;
	assert RAM(30712) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30712))))  severity failure;
	assert RAM(30713) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30713))))  severity failure;
	assert RAM(30714) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(30714))))  severity failure;
	assert RAM(30715) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(30715))))  severity failure;
	assert RAM(30716) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30716))))  severity failure;
	assert RAM(30717) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(30717))))  severity failure;
	assert RAM(30718) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(30718))))  severity failure;
	assert RAM(30719) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(30719))))  severity failure;
	assert RAM(30720) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(30720))))  severity failure;
	assert RAM(30721) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(30721))))  severity failure;
	assert RAM(30722) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(30722))))  severity failure;
	assert RAM(30723) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30723))))  severity failure;
	assert RAM(30724) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(30724))))  severity failure;
	assert RAM(30725) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30725))))  severity failure;
	assert RAM(30726) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(30726))))  severity failure;
	assert RAM(30727) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30727))))  severity failure;
	assert RAM(30728) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(30728))))  severity failure;
	assert RAM(30729) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(30729))))  severity failure;
	assert RAM(30730) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(30730))))  severity failure;
	assert RAM(30731) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(30731))))  severity failure;
	assert RAM(30732) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(30732))))  severity failure;
	assert RAM(30733) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(30733))))  severity failure;
	assert RAM(30734) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(30734))))  severity failure;
	assert RAM(30735) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(30735))))  severity failure;
	assert RAM(30736) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(30736))))  severity failure;
	assert RAM(30737) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30737))))  severity failure;
	assert RAM(30738) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(30738))))  severity failure;
	assert RAM(30739) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(30739))))  severity failure;
	assert RAM(30740) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(30740))))  severity failure;
	assert RAM(30741) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30741))))  severity failure;
	assert RAM(30742) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(30742))))  severity failure;
	assert RAM(30743) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30743))))  severity failure;
	assert RAM(30744) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(30744))))  severity failure;
	assert RAM(30745) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(30745))))  severity failure;
	assert RAM(30746) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(30746))))  severity failure;
	assert RAM(30747) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(30747))))  severity failure;
	assert RAM(30748) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(30748))))  severity failure;
	assert RAM(30749) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(30749))))  severity failure;
	assert RAM(30750) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30750))))  severity failure;
	assert RAM(30751) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(30751))))  severity failure;
	assert RAM(30752) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(30752))))  severity failure;
	assert RAM(30753) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30753))))  severity failure;
	assert RAM(30754) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(30754))))  severity failure;
	assert RAM(30755) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30755))))  severity failure;
	assert RAM(30756) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(30756))))  severity failure;
	assert RAM(30757) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30757))))  severity failure;
	assert RAM(30758) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30758))))  severity failure;
	assert RAM(30759) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30759))))  severity failure;
	assert RAM(30760) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(30760))))  severity failure;
	assert RAM(30761) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30761))))  severity failure;
	assert RAM(30762) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30762))))  severity failure;
	assert RAM(30763) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(30763))))  severity failure;
	assert RAM(30764) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(30764))))  severity failure;
	assert RAM(30765) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(30765))))  severity failure;
	assert RAM(30766) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(30766))))  severity failure;
	assert RAM(30767) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(30767))))  severity failure;
	assert RAM(30768) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(30768))))  severity failure;
	assert RAM(30769) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(30769))))  severity failure;
	assert RAM(30770) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(30770))))  severity failure;
	assert RAM(30771) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(30771))))  severity failure;
	assert RAM(30772) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(30772))))  severity failure;
	assert RAM(30773) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(30773))))  severity failure;
	assert RAM(30774) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(30774))))  severity failure;
	assert RAM(30775) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(30775))))  severity failure;
	assert RAM(30776) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30776))))  severity failure;
	assert RAM(30777) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30777))))  severity failure;
	assert RAM(30778) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(30778))))  severity failure;
	assert RAM(30779) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(30779))))  severity failure;
	assert RAM(30780) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30780))))  severity failure;
	assert RAM(30781) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(30781))))  severity failure;
	assert RAM(30782) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30782))))  severity failure;
	assert RAM(30783) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30783))))  severity failure;
	assert RAM(30784) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(30784))))  severity failure;
	assert RAM(30785) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30785))))  severity failure;
	assert RAM(30786) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30786))))  severity failure;
	assert RAM(30787) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30787))))  severity failure;
	assert RAM(30788) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(30788))))  severity failure;
	assert RAM(30789) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(30789))))  severity failure;
	assert RAM(30790) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(30790))))  severity failure;
	assert RAM(30791) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(30791))))  severity failure;
	assert RAM(30792) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(30792))))  severity failure;
	assert RAM(30793) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(30793))))  severity failure;
	assert RAM(30794) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(30794))))  severity failure;
	assert RAM(30795) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(30795))))  severity failure;
	assert RAM(30796) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(30796))))  severity failure;
	assert RAM(30797) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(30797))))  severity failure;
	assert RAM(30798) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30798))))  severity failure;
	assert RAM(30799) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(30799))))  severity failure;
	assert RAM(30800) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(30800))))  severity failure;
	assert RAM(30801) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(30801))))  severity failure;
	assert RAM(30802) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(30802))))  severity failure;
	assert RAM(30803) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(30803))))  severity failure;
	assert RAM(30804) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30804))))  severity failure;
	assert RAM(30805) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30805))))  severity failure;
	assert RAM(30806) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30806))))  severity failure;
	assert RAM(30807) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(30807))))  severity failure;
	assert RAM(30808) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(30808))))  severity failure;
	assert RAM(30809) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(30809))))  severity failure;
	assert RAM(30810) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(30810))))  severity failure;
	assert RAM(30811) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(30811))))  severity failure;
	assert RAM(30812) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(30812))))  severity failure;
	assert RAM(30813) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(30813))))  severity failure;
	assert RAM(30814) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(30814))))  severity failure;
	assert RAM(30815) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30815))))  severity failure;
	assert RAM(30816) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(30816))))  severity failure;
	assert RAM(30817) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(30817))))  severity failure;
	assert RAM(30818) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(30818))))  severity failure;
	assert RAM(30819) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(30819))))  severity failure;
	assert RAM(30820) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(30820))))  severity failure;
	assert RAM(30821) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(30821))))  severity failure;
	assert RAM(30822) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(30822))))  severity failure;
	assert RAM(30823) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(30823))))  severity failure;
	assert RAM(30824) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(30824))))  severity failure;
	assert RAM(30825) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(30825))))  severity failure;
	assert RAM(30826) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(30826))))  severity failure;
	assert RAM(30827) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(30827))))  severity failure;
	assert RAM(30828) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(30828))))  severity failure;
	assert RAM(30829) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(30829))))  severity failure;
	assert RAM(30830) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(30830))))  severity failure;
	assert RAM(30831) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(30831))))  severity failure;
	assert RAM(30832) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(30832))))  severity failure;
	assert RAM(30833) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30833))))  severity failure;
	assert RAM(30834) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(30834))))  severity failure;
	assert RAM(30835) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(30835))))  severity failure;
	assert RAM(30836) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30836))))  severity failure;
	assert RAM(30837) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(30837))))  severity failure;
	assert RAM(30838) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(30838))))  severity failure;
	assert RAM(30839) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30839))))  severity failure;
	assert RAM(30840) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30840))))  severity failure;
	assert RAM(30841) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30841))))  severity failure;
	assert RAM(30842) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(30842))))  severity failure;
	assert RAM(30843) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(30843))))  severity failure;
	assert RAM(30844) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(30844))))  severity failure;
	assert RAM(30845) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(30845))))  severity failure;
	assert RAM(30846) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(30846))))  severity failure;
	assert RAM(30847) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30847))))  severity failure;
	assert RAM(30848) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(30848))))  severity failure;
	assert RAM(30849) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(30849))))  severity failure;
	assert RAM(30850) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(30850))))  severity failure;
	assert RAM(30851) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30851))))  severity failure;
	assert RAM(30852) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(30852))))  severity failure;
	assert RAM(30853) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(30853))))  severity failure;
	assert RAM(30854) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(30854))))  severity failure;
	assert RAM(30855) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(30855))))  severity failure;
	assert RAM(30856) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(30856))))  severity failure;
	assert RAM(30857) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(30857))))  severity failure;
	assert RAM(30858) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30858))))  severity failure;
	assert RAM(30859) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(30859))))  severity failure;
	assert RAM(30860) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30860))))  severity failure;
	assert RAM(30861) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(30861))))  severity failure;
	assert RAM(30862) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(30862))))  severity failure;
	assert RAM(30863) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(30863))))  severity failure;
	assert RAM(30864) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(30864))))  severity failure;
	assert RAM(30865) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(30865))))  severity failure;
	assert RAM(30866) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(30866))))  severity failure;
	assert RAM(30867) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(30867))))  severity failure;
	assert RAM(30868) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(30868))))  severity failure;
	assert RAM(30869) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(30869))))  severity failure;
	assert RAM(30870) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(30870))))  severity failure;
	assert RAM(30871) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(30871))))  severity failure;
	assert RAM(30872) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(30872))))  severity failure;
	assert RAM(30873) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(30873))))  severity failure;
	assert RAM(30874) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(30874))))  severity failure;
	assert RAM(30875) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(30875))))  severity failure;
	assert RAM(30876) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(30876))))  severity failure;
	assert RAM(30877) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30877))))  severity failure;
	assert RAM(30878) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(30878))))  severity failure;
	assert RAM(30879) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(30879))))  severity failure;
	assert RAM(30880) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30880))))  severity failure;
	assert RAM(30881) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30881))))  severity failure;
	assert RAM(30882) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(30882))))  severity failure;
	assert RAM(30883) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(30883))))  severity failure;
	assert RAM(30884) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(30884))))  severity failure;
	assert RAM(30885) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(30885))))  severity failure;
	assert RAM(30886) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(30886))))  severity failure;
	assert RAM(30887) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(30887))))  severity failure;
	assert RAM(30888) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30888))))  severity failure;
	assert RAM(30889) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(30889))))  severity failure;
	assert RAM(30890) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(30890))))  severity failure;
	assert RAM(30891) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(30891))))  severity failure;
	assert RAM(30892) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(30892))))  severity failure;
	assert RAM(30893) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(30893))))  severity failure;
	assert RAM(30894) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(30894))))  severity failure;
	assert RAM(30895) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30895))))  severity failure;
	assert RAM(30896) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(30896))))  severity failure;
	assert RAM(30897) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30897))))  severity failure;
	assert RAM(30898) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(30898))))  severity failure;
	assert RAM(30899) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30899))))  severity failure;
	assert RAM(30900) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30900))))  severity failure;
	assert RAM(30901) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(30901))))  severity failure;
	assert RAM(30902) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(30902))))  severity failure;
	assert RAM(30903) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(30903))))  severity failure;
	assert RAM(30904) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(30904))))  severity failure;
	assert RAM(30905) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(30905))))  severity failure;
	assert RAM(30906) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(30906))))  severity failure;
	assert RAM(30907) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30907))))  severity failure;
	assert RAM(30908) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(30908))))  severity failure;
	assert RAM(30909) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(30909))))  severity failure;
	assert RAM(30910) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30910))))  severity failure;
	assert RAM(30911) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(30911))))  severity failure;
	assert RAM(30912) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30912))))  severity failure;
	assert RAM(30913) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(30913))))  severity failure;
	assert RAM(30914) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30914))))  severity failure;
	assert RAM(30915) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(30915))))  severity failure;
	assert RAM(30916) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(30916))))  severity failure;
	assert RAM(30917) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30917))))  severity failure;
	assert RAM(30918) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(30918))))  severity failure;
	assert RAM(30919) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(30919))))  severity failure;
	assert RAM(30920) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(30920))))  severity failure;
	assert RAM(30921) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(30921))))  severity failure;
	assert RAM(30922) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(30922))))  severity failure;
	assert RAM(30923) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(30923))))  severity failure;
	assert RAM(30924) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(30924))))  severity failure;
	assert RAM(30925) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(30925))))  severity failure;
	assert RAM(30926) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(30926))))  severity failure;
	assert RAM(30927) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(30927))))  severity failure;
	assert RAM(30928) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(30928))))  severity failure;
	assert RAM(30929) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(30929))))  severity failure;
	assert RAM(30930) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(30930))))  severity failure;
	assert RAM(30931) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(30931))))  severity failure;
	assert RAM(30932) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(30932))))  severity failure;
	assert RAM(30933) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(30933))))  severity failure;
	assert RAM(30934) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(30934))))  severity failure;
	assert RAM(30935) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(30935))))  severity failure;
	assert RAM(30936) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(30936))))  severity failure;
	assert RAM(30937) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(30937))))  severity failure;
	assert RAM(30938) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(30938))))  severity failure;
	assert RAM(30939) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(30939))))  severity failure;
	assert RAM(30940) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30940))))  severity failure;
	assert RAM(30941) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(30941))))  severity failure;
	assert RAM(30942) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(30942))))  severity failure;
	assert RAM(30943) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30943))))  severity failure;
	assert RAM(30944) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(30944))))  severity failure;
	assert RAM(30945) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(30945))))  severity failure;
	assert RAM(30946) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30946))))  severity failure;
	assert RAM(30947) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(30947))))  severity failure;
	assert RAM(30948) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(30948))))  severity failure;
	assert RAM(30949) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(30949))))  severity failure;
	assert RAM(30950) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(30950))))  severity failure;
	assert RAM(30951) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(30951))))  severity failure;
	assert RAM(30952) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(30952))))  severity failure;
	assert RAM(30953) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(30953))))  severity failure;
	assert RAM(30954) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(30954))))  severity failure;
	assert RAM(30955) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(30955))))  severity failure;
	assert RAM(30956) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(30956))))  severity failure;
	assert RAM(30957) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(30957))))  severity failure;
	assert RAM(30958) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(30958))))  severity failure;
	assert RAM(30959) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(30959))))  severity failure;
	assert RAM(30960) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30960))))  severity failure;
	assert RAM(30961) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(30961))))  severity failure;
	assert RAM(30962) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(30962))))  severity failure;
	assert RAM(30963) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(30963))))  severity failure;
	assert RAM(30964) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(30964))))  severity failure;
	assert RAM(30965) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(30965))))  severity failure;
	assert RAM(30966) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(30966))))  severity failure;
	assert RAM(30967) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(30967))))  severity failure;
	assert RAM(30968) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(30968))))  severity failure;
	assert RAM(30969) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(30969))))  severity failure;
	assert RAM(30970) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(30970))))  severity failure;
	assert RAM(30971) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(30971))))  severity failure;
	assert RAM(30972) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(30972))))  severity failure;
	assert RAM(30973) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30973))))  severity failure;
	assert RAM(30974) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(30974))))  severity failure;
	assert RAM(30975) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(30975))))  severity failure;
	assert RAM(30976) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(30976))))  severity failure;
	assert RAM(30977) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(30977))))  severity failure;
	assert RAM(30978) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(30978))))  severity failure;
	assert RAM(30979) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(30979))))  severity failure;
	assert RAM(30980) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(30980))))  severity failure;
	assert RAM(30981) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(30981))))  severity failure;
	assert RAM(30982) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(30982))))  severity failure;
	assert RAM(30983) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(30983))))  severity failure;
	assert RAM(30984) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(30984))))  severity failure;
	assert RAM(30985) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(30985))))  severity failure;
	assert RAM(30986) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(30986))))  severity failure;
	assert RAM(30987) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(30987))))  severity failure;
	assert RAM(30988) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(30988))))  severity failure;
	assert RAM(30989) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(30989))))  severity failure;
	assert RAM(30990) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(30990))))  severity failure;
	assert RAM(30991) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(30991))))  severity failure;
	assert RAM(30992) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(30992))))  severity failure;
	assert RAM(30993) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(30993))))  severity failure;
	assert RAM(30994) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(30994))))  severity failure;
	assert RAM(30995) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(30995))))  severity failure;
	assert RAM(30996) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(30996))))  severity failure;
	assert RAM(30997) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(30997))))  severity failure;
	assert RAM(30998) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(30998))))  severity failure;
	assert RAM(30999) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(30999))))  severity failure;
	assert RAM(31000) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(31000))))  severity failure;
	assert RAM(31001) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(31001))))  severity failure;
	assert RAM(31002) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31002))))  severity failure;
	assert RAM(31003) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(31003))))  severity failure;
	assert RAM(31004) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31004))))  severity failure;
	assert RAM(31005) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31005))))  severity failure;
	assert RAM(31006) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(31006))))  severity failure;
	assert RAM(31007) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(31007))))  severity failure;
	assert RAM(31008) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31008))))  severity failure;
	assert RAM(31009) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(31009))))  severity failure;
	assert RAM(31010) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(31010))))  severity failure;
	assert RAM(31011) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(31011))))  severity failure;
	assert RAM(31012) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(31012))))  severity failure;
	assert RAM(31013) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(31013))))  severity failure;
	assert RAM(31014) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(31014))))  severity failure;
	assert RAM(31015) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31015))))  severity failure;
	assert RAM(31016) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(31016))))  severity failure;
	assert RAM(31017) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31017))))  severity failure;
	assert RAM(31018) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(31018))))  severity failure;
	assert RAM(31019) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(31019))))  severity failure;
	assert RAM(31020) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(31020))))  severity failure;
	assert RAM(31021) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(31021))))  severity failure;
	assert RAM(31022) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(31022))))  severity failure;
	assert RAM(31023) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(31023))))  severity failure;
	assert RAM(31024) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(31024))))  severity failure;
	assert RAM(31025) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31025))))  severity failure;
	assert RAM(31026) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31026))))  severity failure;
	assert RAM(31027) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(31027))))  severity failure;
	assert RAM(31028) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(31028))))  severity failure;
	assert RAM(31029) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31029))))  severity failure;
	assert RAM(31030) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(31030))))  severity failure;
	assert RAM(31031) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(31031))))  severity failure;
	assert RAM(31032) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31032))))  severity failure;
	assert RAM(31033) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(31033))))  severity failure;
	assert RAM(31034) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31034))))  severity failure;
	assert RAM(31035) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31035))))  severity failure;
	assert RAM(31036) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(31036))))  severity failure;
	assert RAM(31037) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(31037))))  severity failure;
	assert RAM(31038) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31038))))  severity failure;
	assert RAM(31039) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(31039))))  severity failure;
	assert RAM(31040) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(31040))))  severity failure;
	assert RAM(31041) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(31041))))  severity failure;
	assert RAM(31042) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31042))))  severity failure;
	assert RAM(31043) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31043))))  severity failure;
	assert RAM(31044) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(31044))))  severity failure;
	assert RAM(31045) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31045))))  severity failure;
	assert RAM(31046) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(31046))))  severity failure;
	assert RAM(31047) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(31047))))  severity failure;
	assert RAM(31048) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31048))))  severity failure;
	assert RAM(31049) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(31049))))  severity failure;
	assert RAM(31050) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(31050))))  severity failure;
	assert RAM(31051) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31051))))  severity failure;
	assert RAM(31052) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31052))))  severity failure;
	assert RAM(31053) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31053))))  severity failure;
	assert RAM(31054) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31054))))  severity failure;
	assert RAM(31055) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31055))))  severity failure;
	assert RAM(31056) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(31056))))  severity failure;
	assert RAM(31057) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31057))))  severity failure;
	assert RAM(31058) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(31058))))  severity failure;
	assert RAM(31059) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(31059))))  severity failure;
	assert RAM(31060) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(31060))))  severity failure;
	assert RAM(31061) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(31061))))  severity failure;
	assert RAM(31062) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(31062))))  severity failure;
	assert RAM(31063) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(31063))))  severity failure;
	assert RAM(31064) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(31064))))  severity failure;
	assert RAM(31065) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31065))))  severity failure;
	assert RAM(31066) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31066))))  severity failure;
	assert RAM(31067) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31067))))  severity failure;
	assert RAM(31068) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(31068))))  severity failure;
	assert RAM(31069) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(31069))))  severity failure;
	assert RAM(31070) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(31070))))  severity failure;
	assert RAM(31071) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31071))))  severity failure;
	assert RAM(31072) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31072))))  severity failure;
	assert RAM(31073) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(31073))))  severity failure;
	assert RAM(31074) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31074))))  severity failure;
	assert RAM(31075) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(31075))))  severity failure;
	assert RAM(31076) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(31076))))  severity failure;
	assert RAM(31077) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31077))))  severity failure;
	assert RAM(31078) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31078))))  severity failure;
	assert RAM(31079) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31079))))  severity failure;
	assert RAM(31080) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31080))))  severity failure;
	assert RAM(31081) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31081))))  severity failure;
	assert RAM(31082) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(31082))))  severity failure;
	assert RAM(31083) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(31083))))  severity failure;
	assert RAM(31084) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(31084))))  severity failure;
	assert RAM(31085) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31085))))  severity failure;
	assert RAM(31086) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(31086))))  severity failure;
	assert RAM(31087) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31087))))  severity failure;
	assert RAM(31088) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(31088))))  severity failure;
	assert RAM(31089) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(31089))))  severity failure;
	assert RAM(31090) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(31090))))  severity failure;
	assert RAM(31091) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31091))))  severity failure;
	assert RAM(31092) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31092))))  severity failure;
	assert RAM(31093) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31093))))  severity failure;
	assert RAM(31094) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(31094))))  severity failure;
	assert RAM(31095) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(31095))))  severity failure;
	assert RAM(31096) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(31096))))  severity failure;
	assert RAM(31097) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31097))))  severity failure;
	assert RAM(31098) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(31098))))  severity failure;
	assert RAM(31099) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(31099))))  severity failure;
	assert RAM(31100) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(31100))))  severity failure;
	assert RAM(31101) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(31101))))  severity failure;
	assert RAM(31102) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(31102))))  severity failure;
	assert RAM(31103) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31103))))  severity failure;
	assert RAM(31104) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(31104))))  severity failure;
	assert RAM(31105) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31105))))  severity failure;
	assert RAM(31106) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(31106))))  severity failure;
	assert RAM(31107) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(31107))))  severity failure;
	assert RAM(31108) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31108))))  severity failure;
	assert RAM(31109) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31109))))  severity failure;
	assert RAM(31110) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(31110))))  severity failure;
	assert RAM(31111) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(31111))))  severity failure;
	assert RAM(31112) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(31112))))  severity failure;
	assert RAM(31113) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(31113))))  severity failure;
	assert RAM(31114) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31114))))  severity failure;
	assert RAM(31115) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(31115))))  severity failure;
	assert RAM(31116) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31116))))  severity failure;
	assert RAM(31117) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(31117))))  severity failure;
	assert RAM(31118) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(31118))))  severity failure;
	assert RAM(31119) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(31119))))  severity failure;
	assert RAM(31120) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(31120))))  severity failure;
	assert RAM(31121) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(31121))))  severity failure;
	assert RAM(31122) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(31122))))  severity failure;
	assert RAM(31123) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(31123))))  severity failure;
	assert RAM(31124) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(31124))))  severity failure;
	assert RAM(31125) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(31125))))  severity failure;
	assert RAM(31126) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(31126))))  severity failure;
	assert RAM(31127) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(31127))))  severity failure;
	assert RAM(31128) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(31128))))  severity failure;
	assert RAM(31129) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(31129))))  severity failure;
	assert RAM(31130) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(31130))))  severity failure;
	assert RAM(31131) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(31131))))  severity failure;
	assert RAM(31132) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31132))))  severity failure;
	assert RAM(31133) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31133))))  severity failure;
	assert RAM(31134) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(31134))))  severity failure;
	assert RAM(31135) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31135))))  severity failure;
	assert RAM(31136) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(31136))))  severity failure;
	assert RAM(31137) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31137))))  severity failure;
	assert RAM(31138) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31138))))  severity failure;
	assert RAM(31139) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(31139))))  severity failure;
	assert RAM(31140) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31140))))  severity failure;
	assert RAM(31141) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(31141))))  severity failure;
	assert RAM(31142) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(31142))))  severity failure;
	assert RAM(31143) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31143))))  severity failure;
	assert RAM(31144) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(31144))))  severity failure;
	assert RAM(31145) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31145))))  severity failure;
	assert RAM(31146) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(31146))))  severity failure;
	assert RAM(31147) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(31147))))  severity failure;
	assert RAM(31148) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(31148))))  severity failure;
	assert RAM(31149) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(31149))))  severity failure;
	assert RAM(31150) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31150))))  severity failure;
	assert RAM(31151) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(31151))))  severity failure;
	assert RAM(31152) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(31152))))  severity failure;
	assert RAM(31153) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(31153))))  severity failure;
	assert RAM(31154) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(31154))))  severity failure;
	assert RAM(31155) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(31155))))  severity failure;
	assert RAM(31156) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(31156))))  severity failure;
	assert RAM(31157) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(31157))))  severity failure;
	assert RAM(31158) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(31158))))  severity failure;
	assert RAM(31159) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(31159))))  severity failure;
	assert RAM(31160) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(31160))))  severity failure;
	assert RAM(31161) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(31161))))  severity failure;
	assert RAM(31162) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(31162))))  severity failure;
	assert RAM(31163) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(31163))))  severity failure;
	assert RAM(31164) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(31164))))  severity failure;
	assert RAM(31165) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(31165))))  severity failure;
	assert RAM(31166) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(31166))))  severity failure;
	assert RAM(31167) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(31167))))  severity failure;
	assert RAM(31168) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(31168))))  severity failure;
	assert RAM(31169) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(31169))))  severity failure;
	assert RAM(31170) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(31170))))  severity failure;
	assert RAM(31171) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31171))))  severity failure;
	assert RAM(31172) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(31172))))  severity failure;
	assert RAM(31173) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(31173))))  severity failure;
	assert RAM(31174) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31174))))  severity failure;
	assert RAM(31175) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(31175))))  severity failure;
	assert RAM(31176) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(31176))))  severity failure;
	assert RAM(31177) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31177))))  severity failure;
	assert RAM(31178) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31178))))  severity failure;
	assert RAM(31179) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31179))))  severity failure;
	assert RAM(31180) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(31180))))  severity failure;
	assert RAM(31181) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(31181))))  severity failure;
	assert RAM(31182) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(31182))))  severity failure;
	assert RAM(31183) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31183))))  severity failure;
	assert RAM(31184) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(31184))))  severity failure;
	assert RAM(31185) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31185))))  severity failure;
	assert RAM(31186) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(31186))))  severity failure;
	assert RAM(31187) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(31187))))  severity failure;
	assert RAM(31188) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(31188))))  severity failure;
	assert RAM(31189) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(31189))))  severity failure;
	assert RAM(31190) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(31190))))  severity failure;
	assert RAM(31191) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31191))))  severity failure;
	assert RAM(31192) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(31192))))  severity failure;
	assert RAM(31193) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(31193))))  severity failure;
	assert RAM(31194) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(31194))))  severity failure;
	assert RAM(31195) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(31195))))  severity failure;
	assert RAM(31196) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31196))))  severity failure;
	assert RAM(31197) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(31197))))  severity failure;
	assert RAM(31198) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(31198))))  severity failure;
	assert RAM(31199) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(31199))))  severity failure;
	assert RAM(31200) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(31200))))  severity failure;
	assert RAM(31201) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(31201))))  severity failure;
	assert RAM(31202) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31202))))  severity failure;
	assert RAM(31203) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(31203))))  severity failure;
	assert RAM(31204) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(31204))))  severity failure;
	assert RAM(31205) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(31205))))  severity failure;
	assert RAM(31206) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(31206))))  severity failure;
	assert RAM(31207) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(31207))))  severity failure;
	assert RAM(31208) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(31208))))  severity failure;
	assert RAM(31209) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(31209))))  severity failure;
	assert RAM(31210) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(31210))))  severity failure;
	assert RAM(31211) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(31211))))  severity failure;
	assert RAM(31212) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(31212))))  severity failure;
	assert RAM(31213) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(31213))))  severity failure;
	assert RAM(31214) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(31214))))  severity failure;
	assert RAM(31215) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31215))))  severity failure;
	assert RAM(31216) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(31216))))  severity failure;
	assert RAM(31217) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(31217))))  severity failure;
	assert RAM(31218) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31218))))  severity failure;
	assert RAM(31219) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(31219))))  severity failure;
	assert RAM(31220) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(31220))))  severity failure;
	assert RAM(31221) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(31221))))  severity failure;
	assert RAM(31222) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(31222))))  severity failure;
	assert RAM(31223) = std_logic_vector(to_unsigned(98,8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(31223))))  severity failure;
	assert RAM(31224) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(31224))))  severity failure;
	assert RAM(31225) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(31225))))  severity failure;
	assert RAM(31226) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(31226))))  severity failure;
	assert RAM(31227) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(31227))))  severity failure;
	assert RAM(31228) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31228))))  severity failure;
	assert RAM(31229) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(31229))))  severity failure;
	assert RAM(31230) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(31230))))  severity failure;
	assert RAM(31231) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31231))))  severity failure;
	assert RAM(31232) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(31232))))  severity failure;
	assert RAM(31233) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(31233))))  severity failure;
	assert RAM(31234) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(31234))))  severity failure;
	assert RAM(31235) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(31235))))  severity failure;
	assert RAM(31236) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31236))))  severity failure;
	assert RAM(31237) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(31237))))  severity failure;
	assert RAM(31238) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(31238))))  severity failure;
	assert RAM(31239) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(31239))))  severity failure;
	assert RAM(31240) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31240))))  severity failure;
	assert RAM(31241) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(31241))))  severity failure;
	assert RAM(31242) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31242))))  severity failure;
	assert RAM(31243) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(31243))))  severity failure;
	assert RAM(31244) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(31244))))  severity failure;
	assert RAM(31245) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31245))))  severity failure;
	assert RAM(31246) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31246))))  severity failure;
	assert RAM(31247) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31247))))  severity failure;
	assert RAM(31248) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(31248))))  severity failure;
	assert RAM(31249) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(31249))))  severity failure;
	assert RAM(31250) = std_logic_vector(to_unsigned(170,8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(31250))))  severity failure;
	assert RAM(31251) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(31251))))  severity failure;
	assert RAM(31252) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(31252))))  severity failure;
	assert RAM(31253) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(31253))))  severity failure;
	assert RAM(31254) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(31254))))  severity failure;
	assert RAM(31255) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31255))))  severity failure;
	assert RAM(31256) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31256))))  severity failure;
	assert RAM(31257) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31257))))  severity failure;
	assert RAM(31258) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31258))))  severity failure;
	assert RAM(31259) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(31259))))  severity failure;
	assert RAM(31260) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31260))))  severity failure;
	assert RAM(31261) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(31261))))  severity failure;
	assert RAM(31262) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(31262))))  severity failure;
	assert RAM(31263) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(31263))))  severity failure;
	assert RAM(31264) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(31264))))  severity failure;
	assert RAM(31265) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(31265))))  severity failure;
	assert RAM(31266) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31266))))  severity failure;
	assert RAM(31267) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(31267))))  severity failure;
	assert RAM(31268) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(31268))))  severity failure;
	assert RAM(31269) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(31269))))  severity failure;
	assert RAM(31270) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(31270))))  severity failure;
	assert RAM(31271) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31271))))  severity failure;
	assert RAM(31272) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(31272))))  severity failure;
	assert RAM(31273) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31273))))  severity failure;
	assert RAM(31274) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(31274))))  severity failure;
	assert RAM(31275) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31275))))  severity failure;
	assert RAM(31276) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31276))))  severity failure;
	assert RAM(31277) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(31277))))  severity failure;
	assert RAM(31278) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(31278))))  severity failure;
	assert RAM(31279) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(31279))))  severity failure;
	assert RAM(31280) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(31280))))  severity failure;
	assert RAM(31281) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(31281))))  severity failure;
	assert RAM(31282) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(31282))))  severity failure;
	assert RAM(31283) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(31283))))  severity failure;
	assert RAM(31284) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(31284))))  severity failure;
	assert RAM(31285) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31285))))  severity failure;
	assert RAM(31286) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(31286))))  severity failure;
	assert RAM(31287) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31287))))  severity failure;
	assert RAM(31288) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(31288))))  severity failure;
	assert RAM(31289) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31289))))  severity failure;
	assert RAM(31290) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(31290))))  severity failure;
	assert RAM(31291) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31291))))  severity failure;
	assert RAM(31292) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(31292))))  severity failure;
	assert RAM(31293) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(31293))))  severity failure;
	assert RAM(31294) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(31294))))  severity failure;
	assert RAM(31295) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(31295))))  severity failure;
	assert RAM(31296) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(31296))))  severity failure;
	assert RAM(31297) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(31297))))  severity failure;
	assert RAM(31298) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(31298))))  severity failure;
	assert RAM(31299) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(31299))))  severity failure;
	assert RAM(31300) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(31300))))  severity failure;
	assert RAM(31301) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(31301))))  severity failure;
	assert RAM(31302) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31302))))  severity failure;
	assert RAM(31303) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(31303))))  severity failure;
	assert RAM(31304) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(31304))))  severity failure;
	assert RAM(31305) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(31305))))  severity failure;
	assert RAM(31306) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31306))))  severity failure;
	assert RAM(31307) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(31307))))  severity failure;
	assert RAM(31308) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(31308))))  severity failure;
	assert RAM(31309) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(31309))))  severity failure;
	assert RAM(31310) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31310))))  severity failure;
	assert RAM(31311) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31311))))  severity failure;
	assert RAM(31312) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31312))))  severity failure;
	assert RAM(31313) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(31313))))  severity failure;
	assert RAM(31314) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(31314))))  severity failure;
	assert RAM(31315) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(31315))))  severity failure;
	assert RAM(31316) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(31316))))  severity failure;
	assert RAM(31317) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(31317))))  severity failure;
	assert RAM(31318) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(31318))))  severity failure;
	assert RAM(31319) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(31319))))  severity failure;
	assert RAM(31320) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31320))))  severity failure;
	assert RAM(31321) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(31321))))  severity failure;
	assert RAM(31322) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(31322))))  severity failure;
	assert RAM(31323) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(31323))))  severity failure;
	assert RAM(31324) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(31324))))  severity failure;
	assert RAM(31325) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(31325))))  severity failure;
	assert RAM(31326) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(31326))))  severity failure;
	assert RAM(31327) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(31327))))  severity failure;
	assert RAM(31328) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(31328))))  severity failure;
	assert RAM(31329) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31329))))  severity failure;
	assert RAM(31330) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(31330))))  severity failure;
	assert RAM(31331) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31331))))  severity failure;
	assert RAM(31332) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(31332))))  severity failure;
	assert RAM(31333) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31333))))  severity failure;
	assert RAM(31334) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(31334))))  severity failure;
	assert RAM(31335) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31335))))  severity failure;
	assert RAM(31336) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31336))))  severity failure;
	assert RAM(31337) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(31337))))  severity failure;
	assert RAM(31338) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31338))))  severity failure;
	assert RAM(31339) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(31339))))  severity failure;
	assert RAM(31340) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(31340))))  severity failure;
	assert RAM(31341) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(31341))))  severity failure;
	assert RAM(31342) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(31342))))  severity failure;
	assert RAM(31343) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31343))))  severity failure;
	assert RAM(31344) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(31344))))  severity failure;
	assert RAM(31345) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(31345))))  severity failure;
	assert RAM(31346) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(31346))))  severity failure;
	assert RAM(31347) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(31347))))  severity failure;
	assert RAM(31348) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31348))))  severity failure;
	assert RAM(31349) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31349))))  severity failure;
	assert RAM(31350) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(31350))))  severity failure;
	assert RAM(31351) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(31351))))  severity failure;
	assert RAM(31352) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(31352))))  severity failure;
	assert RAM(31353) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(31353))))  severity failure;
	assert RAM(31354) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(31354))))  severity failure;
	assert RAM(31355) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31355))))  severity failure;
	assert RAM(31356) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(31356))))  severity failure;
	assert RAM(31357) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(31357))))  severity failure;
	assert RAM(31358) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(31358))))  severity failure;
	assert RAM(31359) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(31359))))  severity failure;
	assert RAM(31360) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31360))))  severity failure;
	assert RAM(31361) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(31361))))  severity failure;
	assert RAM(31362) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(31362))))  severity failure;
	assert RAM(31363) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(31363))))  severity failure;
	assert RAM(31364) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(31364))))  severity failure;
	assert RAM(31365) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31365))))  severity failure;
	assert RAM(31366) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31366))))  severity failure;
	assert RAM(31367) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31367))))  severity failure;
	assert RAM(31368) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31368))))  severity failure;
	assert RAM(31369) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31369))))  severity failure;
	assert RAM(31370) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(31370))))  severity failure;
	assert RAM(31371) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31371))))  severity failure;
	assert RAM(31372) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31372))))  severity failure;
	assert RAM(31373) = std_logic_vector(to_unsigned(204,8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(31373))))  severity failure;
	assert RAM(31374) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31374))))  severity failure;
	assert RAM(31375) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(31375))))  severity failure;
	assert RAM(31376) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(31376))))  severity failure;
	assert RAM(31377) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(31377))))  severity failure;
	assert RAM(31378) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(31378))))  severity failure;
	assert RAM(31379) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31379))))  severity failure;
	assert RAM(31380) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31380))))  severity failure;
	assert RAM(31381) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(31381))))  severity failure;
	assert RAM(31382) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31382))))  severity failure;
	assert RAM(31383) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(31383))))  severity failure;
	assert RAM(31384) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(31384))))  severity failure;
	assert RAM(31385) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(31385))))  severity failure;
	assert RAM(31386) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31386))))  severity failure;
	assert RAM(31387) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(31387))))  severity failure;
	assert RAM(31388) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(31388))))  severity failure;
	assert RAM(31389) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(31389))))  severity failure;
	assert RAM(31390) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(31390))))  severity failure;
	assert RAM(31391) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31391))))  severity failure;
	assert RAM(31392) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(31392))))  severity failure;
	assert RAM(31393) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(31393))))  severity failure;
	assert RAM(31394) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(31394))))  severity failure;
	assert RAM(31395) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31395))))  severity failure;
	assert RAM(31396) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31396))))  severity failure;
	assert RAM(31397) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(31397))))  severity failure;
	assert RAM(31398) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(31398))))  severity failure;
	assert RAM(31399) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(31399))))  severity failure;
	assert RAM(31400) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31400))))  severity failure;
	assert RAM(31401) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31401))))  severity failure;
	assert RAM(31402) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(31402))))  severity failure;
	assert RAM(31403) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(31403))))  severity failure;
	assert RAM(31404) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(31404))))  severity failure;
	assert RAM(31405) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(31405))))  severity failure;
	assert RAM(31406) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31406))))  severity failure;
	assert RAM(31407) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(31407))))  severity failure;
	assert RAM(31408) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(31408))))  severity failure;
	assert RAM(31409) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(31409))))  severity failure;
	assert RAM(31410) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(31410))))  severity failure;
	assert RAM(31411) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(31411))))  severity failure;
	assert RAM(31412) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31412))))  severity failure;
	assert RAM(31413) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(31413))))  severity failure;
	assert RAM(31414) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(31414))))  severity failure;
	assert RAM(31415) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31415))))  severity failure;
	assert RAM(31416) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31416))))  severity failure;
	assert RAM(31417) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(31417))))  severity failure;
	assert RAM(31418) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(31418))))  severity failure;
	assert RAM(31419) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(31419))))  severity failure;
	assert RAM(31420) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31420))))  severity failure;
	assert RAM(31421) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(31421))))  severity failure;
	assert RAM(31422) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31422))))  severity failure;
	assert RAM(31423) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(31423))))  severity failure;
	assert RAM(31424) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(31424))))  severity failure;
	assert RAM(31425) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31425))))  severity failure;
	assert RAM(31426) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(31426))))  severity failure;
	assert RAM(31427) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(31427))))  severity failure;
	assert RAM(31428) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31428))))  severity failure;
	assert RAM(31429) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(31429))))  severity failure;
	assert RAM(31430) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(31430))))  severity failure;
	assert RAM(31431) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(31431))))  severity failure;
	assert RAM(31432) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(31432))))  severity failure;
	assert RAM(31433) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31433))))  severity failure;
	assert RAM(31434) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(31434))))  severity failure;
	assert RAM(31435) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31435))))  severity failure;
	assert RAM(31436) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(31436))))  severity failure;
	assert RAM(31437) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(31437))))  severity failure;
	assert RAM(31438) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31438))))  severity failure;
	assert RAM(31439) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(31439))))  severity failure;
	assert RAM(31440) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31440))))  severity failure;
	assert RAM(31441) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31441))))  severity failure;
	assert RAM(31442) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31442))))  severity failure;
	assert RAM(31443) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(31443))))  severity failure;
	assert RAM(31444) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(31444))))  severity failure;
	assert RAM(31445) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(31445))))  severity failure;
	assert RAM(31446) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(31446))))  severity failure;
	assert RAM(31447) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(31447))))  severity failure;
	assert RAM(31448) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(31448))))  severity failure;
	assert RAM(31449) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(31449))))  severity failure;
	assert RAM(31450) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(31450))))  severity failure;
	assert RAM(31451) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(31451))))  severity failure;
	assert RAM(31452) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(31452))))  severity failure;
	assert RAM(31453) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(31453))))  severity failure;
	assert RAM(31454) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(31454))))  severity failure;
	assert RAM(31455) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31455))))  severity failure;
	assert RAM(31456) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(31456))))  severity failure;
	assert RAM(31457) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(31457))))  severity failure;
	assert RAM(31458) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(31458))))  severity failure;
	assert RAM(31459) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(31459))))  severity failure;
	assert RAM(31460) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(31460))))  severity failure;
	assert RAM(31461) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(31461))))  severity failure;
	assert RAM(31462) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(31462))))  severity failure;
	assert RAM(31463) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31463))))  severity failure;
	assert RAM(31464) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31464))))  severity failure;
	assert RAM(31465) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31465))))  severity failure;
	assert RAM(31466) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(31466))))  severity failure;
	assert RAM(31467) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(31467))))  severity failure;
	assert RAM(31468) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(31468))))  severity failure;
	assert RAM(31469) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(31469))))  severity failure;
	assert RAM(31470) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(31470))))  severity failure;
	assert RAM(31471) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31471))))  severity failure;
	assert RAM(31472) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(31472))))  severity failure;
	assert RAM(31473) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(31473))))  severity failure;
	assert RAM(31474) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(31474))))  severity failure;
	assert RAM(31475) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(31475))))  severity failure;
	assert RAM(31476) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31476))))  severity failure;
	assert RAM(31477) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(31477))))  severity failure;
	assert RAM(31478) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(31478))))  severity failure;
	assert RAM(31479) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(31479))))  severity failure;
	assert RAM(31480) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(31480))))  severity failure;
	assert RAM(31481) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(31481))))  severity failure;
	assert RAM(31482) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(31482))))  severity failure;
	assert RAM(31483) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(31483))))  severity failure;
	assert RAM(31484) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(31484))))  severity failure;
	assert RAM(31485) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(31485))))  severity failure;
	assert RAM(31486) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(31486))))  severity failure;
	assert RAM(31487) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(31487))))  severity failure;
	assert RAM(31488) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(31488))))  severity failure;
	assert RAM(31489) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(31489))))  severity failure;
	assert RAM(31490) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(31490))))  severity failure;
	assert RAM(31491) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(31491))))  severity failure;
	assert RAM(31492) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(31492))))  severity failure;
	assert RAM(31493) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(31493))))  severity failure;
	assert RAM(31494) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(31494))))  severity failure;
	assert RAM(31495) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(31495))))  severity failure;
	assert RAM(31496) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(31496))))  severity failure;
	assert RAM(31497) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(31497))))  severity failure;
	assert RAM(31498) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(31498))))  severity failure;
	assert RAM(31499) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(31499))))  severity failure;
	assert RAM(31500) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(31500))))  severity failure;
	assert RAM(31501) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(31501))))  severity failure;
	assert RAM(31502) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31502))))  severity failure;
	assert RAM(31503) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31503))))  severity failure;
	assert RAM(31504) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(31504))))  severity failure;
	assert RAM(31505) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(31505))))  severity failure;
	assert RAM(31506) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31506))))  severity failure;
	assert RAM(31507) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(31507))))  severity failure;
	assert RAM(31508) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(31508))))  severity failure;
	assert RAM(31509) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(31509))))  severity failure;
	assert RAM(31510) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(31510))))  severity failure;
	assert RAM(31511) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(31511))))  severity failure;
	assert RAM(31512) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(31512))))  severity failure;
	assert RAM(31513) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(31513))))  severity failure;
	assert RAM(31514) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(31514))))  severity failure;
	assert RAM(31515) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(31515))))  severity failure;
	assert RAM(31516) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(31516))))  severity failure;
	assert RAM(31517) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31517))))  severity failure;
	assert RAM(31518) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(31518))))  severity failure;
	assert RAM(31519) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(31519))))  severity failure;
	assert RAM(31520) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(31520))))  severity failure;
	assert RAM(31521) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(31521))))  severity failure;
	assert RAM(31522) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(31522))))  severity failure;
	assert RAM(31523) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(31523))))  severity failure;
	assert RAM(31524) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31524))))  severity failure;
	assert RAM(31525) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(31525))))  severity failure;
	assert RAM(31526) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31526))))  severity failure;
	assert RAM(31527) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31527))))  severity failure;
	assert RAM(31528) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(31528))))  severity failure;
	assert RAM(31529) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31529))))  severity failure;
	assert RAM(31530) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(31530))))  severity failure;
	assert RAM(31531) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(31531))))  severity failure;
	assert RAM(31532) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(31532))))  severity failure;
	assert RAM(31533) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(31533))))  severity failure;
	assert RAM(31534) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(31534))))  severity failure;
	assert RAM(31535) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(31535))))  severity failure;
	assert RAM(31536) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31536))))  severity failure;
	assert RAM(31537) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31537))))  severity failure;
	assert RAM(31538) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31538))))  severity failure;
	assert RAM(31539) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31539))))  severity failure;
	assert RAM(31540) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(31540))))  severity failure;
	assert RAM(31541) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(31541))))  severity failure;
	assert RAM(31542) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(31542))))  severity failure;
	assert RAM(31543) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31543))))  severity failure;
	assert RAM(31544) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(31544))))  severity failure;
	assert RAM(31545) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(31545))))  severity failure;
	assert RAM(31546) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(31546))))  severity failure;
	assert RAM(31547) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(31547))))  severity failure;
	assert RAM(31548) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31548))))  severity failure;
	assert RAM(31549) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(31549))))  severity failure;
	assert RAM(31550) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31550))))  severity failure;
	assert RAM(31551) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(31551))))  severity failure;
	assert RAM(31552) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(31552))))  severity failure;
	assert RAM(31553) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31553))))  severity failure;
	assert RAM(31554) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31554))))  severity failure;
	assert RAM(31555) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(31555))))  severity failure;
	assert RAM(31556) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(31556))))  severity failure;
	assert RAM(31557) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31557))))  severity failure;
	assert RAM(31558) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31558))))  severity failure;
	assert RAM(31559) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(31559))))  severity failure;
	assert RAM(31560) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(31560))))  severity failure;
	assert RAM(31561) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(31561))))  severity failure;
	assert RAM(31562) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(31562))))  severity failure;
	assert RAM(31563) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(31563))))  severity failure;
	assert RAM(31564) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31564))))  severity failure;
	assert RAM(31565) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(31565))))  severity failure;
	assert RAM(31566) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31566))))  severity failure;
	assert RAM(31567) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(31567))))  severity failure;
	assert RAM(31568) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31568))))  severity failure;
	assert RAM(31569) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(31569))))  severity failure;
	assert RAM(31570) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(31570))))  severity failure;
	assert RAM(31571) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(31571))))  severity failure;
	assert RAM(31572) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(31572))))  severity failure;
	assert RAM(31573) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31573))))  severity failure;
	assert RAM(31574) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(31574))))  severity failure;
	assert RAM(31575) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(31575))))  severity failure;
	assert RAM(31576) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(31576))))  severity failure;
	assert RAM(31577) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(31577))))  severity failure;
	assert RAM(31578) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31578))))  severity failure;
	assert RAM(31579) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(31579))))  severity failure;
	assert RAM(31580) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(31580))))  severity failure;
	assert RAM(31581) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(31581))))  severity failure;
	assert RAM(31582) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(31582))))  severity failure;
	assert RAM(31583) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(31583))))  severity failure;
	assert RAM(31584) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(31584))))  severity failure;
	assert RAM(31585) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(31585))))  severity failure;
	assert RAM(31586) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(31586))))  severity failure;
	assert RAM(31587) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(31587))))  severity failure;
	assert RAM(31588) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(31588))))  severity failure;
	assert RAM(31589) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31589))))  severity failure;
	assert RAM(31590) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31590))))  severity failure;
	assert RAM(31591) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(31591))))  severity failure;
	assert RAM(31592) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31592))))  severity failure;
	assert RAM(31593) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(31593))))  severity failure;
	assert RAM(31594) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(31594))))  severity failure;
	assert RAM(31595) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31595))))  severity failure;
	assert RAM(31596) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(31596))))  severity failure;
	assert RAM(31597) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31597))))  severity failure;
	assert RAM(31598) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(31598))))  severity failure;
	assert RAM(31599) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(31599))))  severity failure;
	assert RAM(31600) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(31600))))  severity failure;
	assert RAM(31601) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(31601))))  severity failure;
	assert RAM(31602) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31602))))  severity failure;
	assert RAM(31603) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(31603))))  severity failure;
	assert RAM(31604) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(31604))))  severity failure;
	assert RAM(31605) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(31605))))  severity failure;
	assert RAM(31606) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(31606))))  severity failure;
	assert RAM(31607) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(31607))))  severity failure;
	assert RAM(31608) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31608))))  severity failure;
	assert RAM(31609) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(31609))))  severity failure;
	assert RAM(31610) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(31610))))  severity failure;
	assert RAM(31611) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31611))))  severity failure;
	assert RAM(31612) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(31612))))  severity failure;
	assert RAM(31613) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31613))))  severity failure;
	assert RAM(31614) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(31614))))  severity failure;
	assert RAM(31615) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(31615))))  severity failure;
	assert RAM(31616) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31616))))  severity failure;
	assert RAM(31617) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(31617))))  severity failure;
	assert RAM(31618) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31618))))  severity failure;
	assert RAM(31619) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31619))))  severity failure;
	assert RAM(31620) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(31620))))  severity failure;
	assert RAM(31621) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(31621))))  severity failure;
	assert RAM(31622) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31622))))  severity failure;
	assert RAM(31623) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31623))))  severity failure;
	assert RAM(31624) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31624))))  severity failure;
	assert RAM(31625) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(31625))))  severity failure;
	assert RAM(31626) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(31626))))  severity failure;
	assert RAM(31627) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(31627))))  severity failure;
	assert RAM(31628) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(31628))))  severity failure;
	assert RAM(31629) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31629))))  severity failure;
	assert RAM(31630) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(31630))))  severity failure;
	assert RAM(31631) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31631))))  severity failure;
	assert RAM(31632) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(31632))))  severity failure;
	assert RAM(31633) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(31633))))  severity failure;
	assert RAM(31634) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(31634))))  severity failure;
	assert RAM(31635) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31635))))  severity failure;
	assert RAM(31636) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(31636))))  severity failure;
	assert RAM(31637) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(31637))))  severity failure;
	assert RAM(31638) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(31638))))  severity failure;
	assert RAM(31639) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(31639))))  severity failure;
	assert RAM(31640) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31640))))  severity failure;
	assert RAM(31641) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31641))))  severity failure;
	assert RAM(31642) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(31642))))  severity failure;
	assert RAM(31643) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(31643))))  severity failure;
	assert RAM(31644) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(31644))))  severity failure;
	assert RAM(31645) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31645))))  severity failure;
	assert RAM(31646) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(31646))))  severity failure;
	assert RAM(31647) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(31647))))  severity failure;
	assert RAM(31648) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(31648))))  severity failure;
	assert RAM(31649) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(31649))))  severity failure;
	assert RAM(31650) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31650))))  severity failure;
	assert RAM(31651) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31651))))  severity failure;
	assert RAM(31652) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(31652))))  severity failure;
	assert RAM(31653) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(31653))))  severity failure;
	assert RAM(31654) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31654))))  severity failure;
	assert RAM(31655) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(31655))))  severity failure;
	assert RAM(31656) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31656))))  severity failure;
	assert RAM(31657) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31657))))  severity failure;
	assert RAM(31658) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31658))))  severity failure;
	assert RAM(31659) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(31659))))  severity failure;
	assert RAM(31660) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31660))))  severity failure;
	assert RAM(31661) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(31661))))  severity failure;
	assert RAM(31662) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31662))))  severity failure;
	assert RAM(31663) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31663))))  severity failure;
	assert RAM(31664) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(31664))))  severity failure;
	assert RAM(31665) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(31665))))  severity failure;
	assert RAM(31666) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(31666))))  severity failure;
	assert RAM(31667) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(31667))))  severity failure;
	assert RAM(31668) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(31668))))  severity failure;
	assert RAM(31669) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(31669))))  severity failure;
	assert RAM(31670) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(31670))))  severity failure;
	assert RAM(31671) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31671))))  severity failure;
	assert RAM(31672) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(31672))))  severity failure;
	assert RAM(31673) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(31673))))  severity failure;
	assert RAM(31674) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31674))))  severity failure;
	assert RAM(31675) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(31675))))  severity failure;
	assert RAM(31676) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31676))))  severity failure;
	assert RAM(31677) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(31677))))  severity failure;
	assert RAM(31678) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(31678))))  severity failure;
	assert RAM(31679) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(31679))))  severity failure;
	assert RAM(31680) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(31680))))  severity failure;
	assert RAM(31681) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(31681))))  severity failure;
	assert RAM(31682) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31682))))  severity failure;
	assert RAM(31683) = std_logic_vector(to_unsigned(56,8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(31683))))  severity failure;
	assert RAM(31684) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(31684))))  severity failure;
	assert RAM(31685) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31685))))  severity failure;
	assert RAM(31686) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31686))))  severity failure;
	assert RAM(31687) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(31687))))  severity failure;
	assert RAM(31688) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(31688))))  severity failure;
	assert RAM(31689) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31689))))  severity failure;
	assert RAM(31690) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(31690))))  severity failure;
	assert RAM(31691) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(31691))))  severity failure;
	assert RAM(31692) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(31692))))  severity failure;
	assert RAM(31693) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(31693))))  severity failure;
	assert RAM(31694) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(31694))))  severity failure;
	assert RAM(31695) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(31695))))  severity failure;
	assert RAM(31696) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(31696))))  severity failure;
	assert RAM(31697) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(31697))))  severity failure;
	assert RAM(31698) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(31698))))  severity failure;
	assert RAM(31699) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(31699))))  severity failure;
	assert RAM(31700) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(31700))))  severity failure;
	assert RAM(31701) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(31701))))  severity failure;
	assert RAM(31702) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(31702))))  severity failure;
	assert RAM(31703) = std_logic_vector(to_unsigned(5,8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(31703))))  severity failure;
	assert RAM(31704) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31704))))  severity failure;
	assert RAM(31705) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(31705))))  severity failure;
	assert RAM(31706) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31706))))  severity failure;
	assert RAM(31707) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(31707))))  severity failure;
	assert RAM(31708) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(31708))))  severity failure;
	assert RAM(31709) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31709))))  severity failure;
	assert RAM(31710) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(31710))))  severity failure;
	assert RAM(31711) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(31711))))  severity failure;
	assert RAM(31712) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(31712))))  severity failure;
	assert RAM(31713) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(31713))))  severity failure;
	assert RAM(31714) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(31714))))  severity failure;
	assert RAM(31715) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(31715))))  severity failure;
	assert RAM(31716) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(31716))))  severity failure;
	assert RAM(31717) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31717))))  severity failure;
	assert RAM(31718) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31718))))  severity failure;
	assert RAM(31719) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(31719))))  severity failure;
	assert RAM(31720) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(31720))))  severity failure;
	assert RAM(31721) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(31721))))  severity failure;
	assert RAM(31722) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31722))))  severity failure;
	assert RAM(31723) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(31723))))  severity failure;
	assert RAM(31724) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(31724))))  severity failure;
	assert RAM(31725) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31725))))  severity failure;
	assert RAM(31726) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(31726))))  severity failure;
	assert RAM(31727) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(31727))))  severity failure;
	assert RAM(31728) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(31728))))  severity failure;
	assert RAM(31729) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(31729))))  severity failure;
	assert RAM(31730) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(31730))))  severity failure;
	assert RAM(31731) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(31731))))  severity failure;
	assert RAM(31732) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(31732))))  severity failure;
	assert RAM(31733) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(31733))))  severity failure;
	assert RAM(31734) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31734))))  severity failure;
	assert RAM(31735) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(31735))))  severity failure;
	assert RAM(31736) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(31736))))  severity failure;
	assert RAM(31737) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31737))))  severity failure;
	assert RAM(31738) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(31738))))  severity failure;
	assert RAM(31739) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(31739))))  severity failure;
	assert RAM(31740) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(31740))))  severity failure;
	assert RAM(31741) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(31741))))  severity failure;
	assert RAM(31742) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(31742))))  severity failure;
	assert RAM(31743) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(31743))))  severity failure;
	assert RAM(31744) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(31744))))  severity failure;
	assert RAM(31745) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31745))))  severity failure;
	assert RAM(31746) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(31746))))  severity failure;
	assert RAM(31747) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(31747))))  severity failure;
	assert RAM(31748) = std_logic_vector(to_unsigned(198,8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(31748))))  severity failure;
	assert RAM(31749) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(31749))))  severity failure;
	assert RAM(31750) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(31750))))  severity failure;
	assert RAM(31751) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(31751))))  severity failure;
	assert RAM(31752) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31752))))  severity failure;
	assert RAM(31753) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(31753))))  severity failure;
	assert RAM(31754) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(31754))))  severity failure;
	assert RAM(31755) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(31755))))  severity failure;
	assert RAM(31756) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(31756))))  severity failure;
	assert RAM(31757) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(31757))))  severity failure;
	assert RAM(31758) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(31758))))  severity failure;
	assert RAM(31759) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(31759))))  severity failure;
	assert RAM(31760) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(31760))))  severity failure;
	assert RAM(31761) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31761))))  severity failure;
	assert RAM(31762) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31762))))  severity failure;
	assert RAM(31763) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31763))))  severity failure;
	assert RAM(31764) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(31764))))  severity failure;
	assert RAM(31765) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(31765))))  severity failure;
	assert RAM(31766) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(31766))))  severity failure;
	assert RAM(31767) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(31767))))  severity failure;
	assert RAM(31768) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(31768))))  severity failure;
	assert RAM(31769) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(31769))))  severity failure;
	assert RAM(31770) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(31770))))  severity failure;
	assert RAM(31771) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(31771))))  severity failure;
	assert RAM(31772) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(31772))))  severity failure;
	assert RAM(31773) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(31773))))  severity failure;
	assert RAM(31774) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31774))))  severity failure;
	assert RAM(31775) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(31775))))  severity failure;
	assert RAM(31776) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(31776))))  severity failure;
	assert RAM(31777) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(31777))))  severity failure;
	assert RAM(31778) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(31778))))  severity failure;
	assert RAM(31779) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(31779))))  severity failure;
	assert RAM(31780) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(31780))))  severity failure;
	assert RAM(31781) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(31781))))  severity failure;
	assert RAM(31782) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31782))))  severity failure;
	assert RAM(31783) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(31783))))  severity failure;
	assert RAM(31784) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(31784))))  severity failure;
	assert RAM(31785) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(31785))))  severity failure;
	assert RAM(31786) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(31786))))  severity failure;
	assert RAM(31787) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(31787))))  severity failure;
	assert RAM(31788) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(31788))))  severity failure;
	assert RAM(31789) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(31789))))  severity failure;
	assert RAM(31790) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(31790))))  severity failure;
	assert RAM(31791) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31791))))  severity failure;
	assert RAM(31792) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31792))))  severity failure;
	assert RAM(31793) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(31793))))  severity failure;
	assert RAM(31794) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31794))))  severity failure;
	assert RAM(31795) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(31795))))  severity failure;
	assert RAM(31796) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(31796))))  severity failure;
	assert RAM(31797) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(31797))))  severity failure;
	assert RAM(31798) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31798))))  severity failure;
	assert RAM(31799) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31799))))  severity failure;
	assert RAM(31800) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(31800))))  severity failure;
	assert RAM(31801) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(31801))))  severity failure;
	assert RAM(31802) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31802))))  severity failure;
	assert RAM(31803) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(31803))))  severity failure;
	assert RAM(31804) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31804))))  severity failure;
	assert RAM(31805) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(31805))))  severity failure;
	assert RAM(31806) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(31806))))  severity failure;
	assert RAM(31807) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(31807))))  severity failure;
	assert RAM(31808) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(31808))))  severity failure;
	assert RAM(31809) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(31809))))  severity failure;
	assert RAM(31810) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31810))))  severity failure;
	assert RAM(31811) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(31811))))  severity failure;
	assert RAM(31812) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(31812))))  severity failure;
	assert RAM(31813) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31813))))  severity failure;
	assert RAM(31814) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31814))))  severity failure;
	assert RAM(31815) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31815))))  severity failure;
	assert RAM(31816) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(31816))))  severity failure;
	assert RAM(31817) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(31817))))  severity failure;
	assert RAM(31818) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(31818))))  severity failure;
	assert RAM(31819) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31819))))  severity failure;
	assert RAM(31820) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(31820))))  severity failure;
	assert RAM(31821) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31821))))  severity failure;
	assert RAM(31822) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(31822))))  severity failure;
	assert RAM(31823) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(31823))))  severity failure;
	assert RAM(31824) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(31824))))  severity failure;
	assert RAM(31825) = std_logic_vector(to_unsigned(153,8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(31825))))  severity failure;
	assert RAM(31826) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(31826))))  severity failure;
	assert RAM(31827) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(31827))))  severity failure;
	assert RAM(31828) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31828))))  severity failure;
	assert RAM(31829) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(31829))))  severity failure;
	assert RAM(31830) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(31830))))  severity failure;
	assert RAM(31831) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(31831))))  severity failure;
	assert RAM(31832) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(31832))))  severity failure;
	assert RAM(31833) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(31833))))  severity failure;
	assert RAM(31834) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(31834))))  severity failure;
	assert RAM(31835) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(31835))))  severity failure;
	assert RAM(31836) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(31836))))  severity failure;
	assert RAM(31837) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(31837))))  severity failure;
	assert RAM(31838) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(31838))))  severity failure;
	assert RAM(31839) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31839))))  severity failure;
	assert RAM(31840) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(31840))))  severity failure;
	assert RAM(31841) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(31841))))  severity failure;
	assert RAM(31842) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(31842))))  severity failure;
	assert RAM(31843) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(31843))))  severity failure;
	assert RAM(31844) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(31844))))  severity failure;
	assert RAM(31845) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31845))))  severity failure;
	assert RAM(31846) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(31846))))  severity failure;
	assert RAM(31847) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31847))))  severity failure;
	assert RAM(31848) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31848))))  severity failure;
	assert RAM(31849) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(31849))))  severity failure;
	assert RAM(31850) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(31850))))  severity failure;
	assert RAM(31851) = std_logic_vector(to_unsigned(254,8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(31851))))  severity failure;
	assert RAM(31852) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(31852))))  severity failure;
	assert RAM(31853) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(31853))))  severity failure;
	assert RAM(31854) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(31854))))  severity failure;
	assert RAM(31855) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(31855))))  severity failure;
	assert RAM(31856) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(31856))))  severity failure;
	assert RAM(31857) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(31857))))  severity failure;
	assert RAM(31858) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(31858))))  severity failure;
	assert RAM(31859) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(31859))))  severity failure;
	assert RAM(31860) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(31860))))  severity failure;
	assert RAM(31861) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(31861))))  severity failure;
	assert RAM(31862) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(31862))))  severity failure;
	assert RAM(31863) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(31863))))  severity failure;
	assert RAM(31864) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(31864))))  severity failure;
	assert RAM(31865) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(31865))))  severity failure;
	assert RAM(31866) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(31866))))  severity failure;
	assert RAM(31867) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(31867))))  severity failure;
	assert RAM(31868) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31868))))  severity failure;
	assert RAM(31869) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(31869))))  severity failure;
	assert RAM(31870) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(31870))))  severity failure;
	assert RAM(31871) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(31871))))  severity failure;
	assert RAM(31872) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(31872))))  severity failure;
	assert RAM(31873) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31873))))  severity failure;
	assert RAM(31874) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(31874))))  severity failure;
	assert RAM(31875) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(31875))))  severity failure;
	assert RAM(31876) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(31876))))  severity failure;
	assert RAM(31877) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(31877))))  severity failure;
	assert RAM(31878) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(31878))))  severity failure;
	assert RAM(31879) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(31879))))  severity failure;
	assert RAM(31880) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31880))))  severity failure;
	assert RAM(31881) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31881))))  severity failure;
	assert RAM(31882) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(31882))))  severity failure;
	assert RAM(31883) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(31883))))  severity failure;
	assert RAM(31884) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(31884))))  severity failure;
	assert RAM(31885) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(31885))))  severity failure;
	assert RAM(31886) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(31886))))  severity failure;
	assert RAM(31887) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(31887))))  severity failure;
	assert RAM(31888) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(31888))))  severity failure;
	assert RAM(31889) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(31889))))  severity failure;
	assert RAM(31890) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(31890))))  severity failure;
	assert RAM(31891) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(31891))))  severity failure;
	assert RAM(31892) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(31892))))  severity failure;
	assert RAM(31893) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(31893))))  severity failure;
	assert RAM(31894) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(31894))))  severity failure;
	assert RAM(31895) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(31895))))  severity failure;
	assert RAM(31896) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(31896))))  severity failure;
	assert RAM(31897) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(31897))))  severity failure;
	assert RAM(31898) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(31898))))  severity failure;
	assert RAM(31899) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(31899))))  severity failure;
	assert RAM(31900) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(31900))))  severity failure;
	assert RAM(31901) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31901))))  severity failure;
	assert RAM(31902) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(31902))))  severity failure;
	assert RAM(31903) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(31903))))  severity failure;
	assert RAM(31904) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(31904))))  severity failure;
	assert RAM(31905) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31905))))  severity failure;
	assert RAM(31906) = std_logic_vector(to_unsigned(184,8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(31906))))  severity failure;
	assert RAM(31907) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(31907))))  severity failure;
	assert RAM(31908) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31908))))  severity failure;
	assert RAM(31909) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(31909))))  severity failure;
	assert RAM(31910) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(31910))))  severity failure;
	assert RAM(31911) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31911))))  severity failure;
	assert RAM(31912) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(31912))))  severity failure;
	assert RAM(31913) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31913))))  severity failure;
	assert RAM(31914) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(31914))))  severity failure;
	assert RAM(31915) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(31915))))  severity failure;
	assert RAM(31916) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(31916))))  severity failure;
	assert RAM(31917) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(31917))))  severity failure;
	assert RAM(31918) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(31918))))  severity failure;
	assert RAM(31919) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(31919))))  severity failure;
	assert RAM(31920) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(31920))))  severity failure;
	assert RAM(31921) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31921))))  severity failure;
	assert RAM(31922) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(31922))))  severity failure;
	assert RAM(31923) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(31923))))  severity failure;
	assert RAM(31924) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(31924))))  severity failure;
	assert RAM(31925) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(31925))))  severity failure;
	assert RAM(31926) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(31926))))  severity failure;
	assert RAM(31927) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(31927))))  severity failure;
	assert RAM(31928) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(31928))))  severity failure;
	assert RAM(31929) = std_logic_vector(to_unsigned(155,8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(31929))))  severity failure;
	assert RAM(31930) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(31930))))  severity failure;
	assert RAM(31931) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(31931))))  severity failure;
	assert RAM(31932) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(31932))))  severity failure;
	assert RAM(31933) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(31933))))  severity failure;
	assert RAM(31934) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(31934))))  severity failure;
	assert RAM(31935) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(31935))))  severity failure;
	assert RAM(31936) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31936))))  severity failure;
	assert RAM(31937) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(31937))))  severity failure;
	assert RAM(31938) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(31938))))  severity failure;
	assert RAM(31939) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(31939))))  severity failure;
	assert RAM(31940) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(31940))))  severity failure;
	assert RAM(31941) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31941))))  severity failure;
	assert RAM(31942) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(31942))))  severity failure;
	assert RAM(31943) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(31943))))  severity failure;
	assert RAM(31944) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(31944))))  severity failure;
	assert RAM(31945) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(31945))))  severity failure;
	assert RAM(31946) = std_logic_vector(to_unsigned(158,8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(31946))))  severity failure;
	assert RAM(31947) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(31947))))  severity failure;
	assert RAM(31948) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(31948))))  severity failure;
	assert RAM(31949) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(31949))))  severity failure;
	assert RAM(31950) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(31950))))  severity failure;
	assert RAM(31951) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(31951))))  severity failure;
	assert RAM(31952) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(31952))))  severity failure;
	assert RAM(31953) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(31953))))  severity failure;
	assert RAM(31954) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(31954))))  severity failure;
	assert RAM(31955) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(31955))))  severity failure;
	assert RAM(31956) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(31956))))  severity failure;
	assert RAM(31957) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31957))))  severity failure;
	assert RAM(31958) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(31958))))  severity failure;
	assert RAM(31959) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(31959))))  severity failure;
	assert RAM(31960) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(31960))))  severity failure;
	assert RAM(31961) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(31961))))  severity failure;
	assert RAM(31962) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(31962))))  severity failure;
	assert RAM(31963) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(31963))))  severity failure;
	assert RAM(31964) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(31964))))  severity failure;
	assert RAM(31965) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(31965))))  severity failure;
	assert RAM(31966) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(31966))))  severity failure;
	assert RAM(31967) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(31967))))  severity failure;
	assert RAM(31968) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(31968))))  severity failure;
	assert RAM(31969) = std_logic_vector(to_unsigned(3,8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(31969))))  severity failure;
	assert RAM(31970) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(31970))))  severity failure;
	assert RAM(31971) = std_logic_vector(to_unsigned(88,8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(31971))))  severity failure;
	assert RAM(31972) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(31972))))  severity failure;
	assert RAM(31973) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(31973))))  severity failure;
	assert RAM(31974) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(31974))))  severity failure;
	assert RAM(31975) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(31975))))  severity failure;
	assert RAM(31976) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(31976))))  severity failure;
	assert RAM(31977) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(31977))))  severity failure;
	assert RAM(31978) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31978))))  severity failure;
	assert RAM(31979) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(31979))))  severity failure;
	assert RAM(31980) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(31980))))  severity failure;
	assert RAM(31981) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(31981))))  severity failure;
	assert RAM(31982) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(31982))))  severity failure;
	assert RAM(31983) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(31983))))  severity failure;
	assert RAM(31984) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(31984))))  severity failure;
	assert RAM(31985) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(31985))))  severity failure;
	assert RAM(31986) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(31986))))  severity failure;
	assert RAM(31987) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(31987))))  severity failure;
	assert RAM(31988) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(31988))))  severity failure;
	assert RAM(31989) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(31989))))  severity failure;
	assert RAM(31990) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(31990))))  severity failure;
	assert RAM(31991) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(31991))))  severity failure;
	assert RAM(31992) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(31992))))  severity failure;
	assert RAM(31993) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(31993))))  severity failure;
	assert RAM(31994) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(31994))))  severity failure;
	assert RAM(31995) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(31995))))  severity failure;
	assert RAM(31996) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(31996))))  severity failure;
	assert RAM(31997) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(31997))))  severity failure;
	assert RAM(31998) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(31998))))  severity failure;
	assert RAM(31999) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(31999))))  severity failure;
	assert RAM(32000) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(32000))))  severity failure;
	assert RAM(32001) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(32001))))  severity failure;
	assert RAM(32002) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32002))))  severity failure;
	assert RAM(32003) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(32003))))  severity failure;
	assert RAM(32004) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(32004))))  severity failure;
	assert RAM(32005) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(32005))))  severity failure;
	assert RAM(32006) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(32006))))  severity failure;
	assert RAM(32007) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(32007))))  severity failure;
	assert RAM(32008) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32008))))  severity failure;
	assert RAM(32009) = std_logic_vector(to_unsigned(240,8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(32009))))  severity failure;
	assert RAM(32010) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(32010))))  severity failure;
	assert RAM(32011) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(32011))))  severity failure;
	assert RAM(32012) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(32012))))  severity failure;
	assert RAM(32013) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(32013))))  severity failure;
	assert RAM(32014) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(32014))))  severity failure;
	assert RAM(32015) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(32015))))  severity failure;
	assert RAM(32016) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32016))))  severity failure;
	assert RAM(32017) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(32017))))  severity failure;
	assert RAM(32018) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32018))))  severity failure;
	assert RAM(32019) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(32019))))  severity failure;
	assert RAM(32020) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(32020))))  severity failure;
	assert RAM(32021) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(32021))))  severity failure;
	assert RAM(32022) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(32022))))  severity failure;
	assert RAM(32023) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32023))))  severity failure;
	assert RAM(32024) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(32024))))  severity failure;
	assert RAM(32025) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(32025))))  severity failure;
	assert RAM(32026) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(32026))))  severity failure;
	assert RAM(32027) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(32027))))  severity failure;
	assert RAM(32028) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(32028))))  severity failure;
	assert RAM(32029) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(32029))))  severity failure;
	assert RAM(32030) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(32030))))  severity failure;
	assert RAM(32031) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32031))))  severity failure;
	assert RAM(32032) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(32032))))  severity failure;
	assert RAM(32033) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(32033))))  severity failure;
	assert RAM(32034) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(32034))))  severity failure;
	assert RAM(32035) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(32035))))  severity failure;
	assert RAM(32036) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(32036))))  severity failure;
	assert RAM(32037) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(32037))))  severity failure;
	assert RAM(32038) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(32038))))  severity failure;
	assert RAM(32039) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(32039))))  severity failure;
	assert RAM(32040) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(32040))))  severity failure;
	assert RAM(32041) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(32041))))  severity failure;
	assert RAM(32042) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(32042))))  severity failure;
	assert RAM(32043) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32043))))  severity failure;
	assert RAM(32044) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32044))))  severity failure;
	assert RAM(32045) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(32045))))  severity failure;
	assert RAM(32046) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(32046))))  severity failure;
	assert RAM(32047) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(32047))))  severity failure;
	assert RAM(32048) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32048))))  severity failure;
	assert RAM(32049) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32049))))  severity failure;
	assert RAM(32050) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(32050))))  severity failure;
	assert RAM(32051) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(32051))))  severity failure;
	assert RAM(32052) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(32052))))  severity failure;
	assert RAM(32053) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(32053))))  severity failure;
	assert RAM(32054) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(32054))))  severity failure;
	assert RAM(32055) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(32055))))  severity failure;
	assert RAM(32056) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(32056))))  severity failure;
	assert RAM(32057) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(32057))))  severity failure;
	assert RAM(32058) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(32058))))  severity failure;
	assert RAM(32059) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(32059))))  severity failure;
	assert RAM(32060) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(32060))))  severity failure;
	assert RAM(32061) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32061))))  severity failure;
	assert RAM(32062) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32062))))  severity failure;
	assert RAM(32063) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(32063))))  severity failure;
	assert RAM(32064) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(32064))))  severity failure;
	assert RAM(32065) = std_logic_vector(to_unsigned(77,8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(32065))))  severity failure;
	assert RAM(32066) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(32066))))  severity failure;
	assert RAM(32067) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(32067))))  severity failure;
	assert RAM(32068) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(32068))))  severity failure;
	assert RAM(32069) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(32069))))  severity failure;
	assert RAM(32070) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(32070))))  severity failure;
	assert RAM(32071) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32071))))  severity failure;
	assert RAM(32072) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(32072))))  severity failure;
	assert RAM(32073) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(32073))))  severity failure;
	assert RAM(32074) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32074))))  severity failure;
	assert RAM(32075) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(32075))))  severity failure;
	assert RAM(32076) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(32076))))  severity failure;
	assert RAM(32077) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(32077))))  severity failure;
	assert RAM(32078) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32078))))  severity failure;
	assert RAM(32079) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(32079))))  severity failure;
	assert RAM(32080) = std_logic_vector(to_unsigned(62,8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(32080))))  severity failure;
	assert RAM(32081) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(32081))))  severity failure;
	assert RAM(32082) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32082))))  severity failure;
	assert RAM(32083) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32083))))  severity failure;
	assert RAM(32084) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(32084))))  severity failure;
	assert RAM(32085) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(32085))))  severity failure;
	assert RAM(32086) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(32086))))  severity failure;
	assert RAM(32087) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(32087))))  severity failure;
	assert RAM(32088) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(32088))))  severity failure;
	assert RAM(32089) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(32089))))  severity failure;
	assert RAM(32090) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(32090))))  severity failure;
	assert RAM(32091) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(32091))))  severity failure;
	assert RAM(32092) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32092))))  severity failure;
	assert RAM(32093) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(32093))))  severity failure;
	assert RAM(32094) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(32094))))  severity failure;
	assert RAM(32095) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(32095))))  severity failure;
	assert RAM(32096) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32096))))  severity failure;
	assert RAM(32097) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(32097))))  severity failure;
	assert RAM(32098) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(32098))))  severity failure;
	assert RAM(32099) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(32099))))  severity failure;
	assert RAM(32100) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(32100))))  severity failure;
	assert RAM(32101) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(32101))))  severity failure;
	assert RAM(32102) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32102))))  severity failure;
	assert RAM(32103) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(32103))))  severity failure;
	assert RAM(32104) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(32104))))  severity failure;
	assert RAM(32105) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(32105))))  severity failure;
	assert RAM(32106) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(32106))))  severity failure;
	assert RAM(32107) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(32107))))  severity failure;
	assert RAM(32108) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(32108))))  severity failure;
	assert RAM(32109) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(32109))))  severity failure;
	assert RAM(32110) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(32110))))  severity failure;
	assert RAM(32111) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(32111))))  severity failure;
	assert RAM(32112) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(32112))))  severity failure;
	assert RAM(32113) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(32113))))  severity failure;
	assert RAM(32114) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(32114))))  severity failure;
	assert RAM(32115) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(32115))))  severity failure;
	assert RAM(32116) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(32116))))  severity failure;
	assert RAM(32117) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(32117))))  severity failure;
	assert RAM(32118) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(32118))))  severity failure;
	assert RAM(32119) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(32119))))  severity failure;
	assert RAM(32120) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(32120))))  severity failure;
	assert RAM(32121) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(32121))))  severity failure;
	assert RAM(32122) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(32122))))  severity failure;
	assert RAM(32123) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(32123))))  severity failure;
	assert RAM(32124) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(32124))))  severity failure;
	assert RAM(32125) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(32125))))  severity failure;
	assert RAM(32126) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(32126))))  severity failure;
	assert RAM(32127) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(32127))))  severity failure;
	assert RAM(32128) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(32128))))  severity failure;
	assert RAM(32129) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(32129))))  severity failure;
	assert RAM(32130) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32130))))  severity failure;
	assert RAM(32131) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(32131))))  severity failure;
	assert RAM(32132) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32132))))  severity failure;
	assert RAM(32133) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(32133))))  severity failure;
	assert RAM(32134) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(32134))))  severity failure;
	assert RAM(32135) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(32135))))  severity failure;
	assert RAM(32136) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(32136))))  severity failure;
	assert RAM(32137) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(32137))))  severity failure;
	assert RAM(32138) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(32138))))  severity failure;
	assert RAM(32139) = std_logic_vector(to_unsigned(115,8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(32139))))  severity failure;
	assert RAM(32140) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(32140))))  severity failure;
	assert RAM(32141) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(32141))))  severity failure;
	assert RAM(32142) = std_logic_vector(to_unsigned(200,8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(32142))))  severity failure;
	assert RAM(32143) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(32143))))  severity failure;
	assert RAM(32144) = std_logic_vector(to_unsigned(25,8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(32144))))  severity failure;
	assert RAM(32145) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32145))))  severity failure;
	assert RAM(32146) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(32146))))  severity failure;
	assert RAM(32147) = std_logic_vector(to_unsigned(125,8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(32147))))  severity failure;
	assert RAM(32148) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(32148))))  severity failure;
	assert RAM(32149) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(32149))))  severity failure;
	assert RAM(32150) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(32150))))  severity failure;
	assert RAM(32151) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(32151))))  severity failure;
	assert RAM(32152) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(32152))))  severity failure;
	assert RAM(32153) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(32153))))  severity failure;
	assert RAM(32154) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(32154))))  severity failure;
	assert RAM(32155) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(32155))))  severity failure;
	assert RAM(32156) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32156))))  severity failure;
	assert RAM(32157) = std_logic_vector(to_unsigned(14,8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(32157))))  severity failure;
	assert RAM(32158) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32158))))  severity failure;
	assert RAM(32159) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(32159))))  severity failure;
	assert RAM(32160) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(32160))))  severity failure;
	assert RAM(32161) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(32161))))  severity failure;
	assert RAM(32162) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(32162))))  severity failure;
	assert RAM(32163) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(32163))))  severity failure;
	assert RAM(32164) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(32164))))  severity failure;
	assert RAM(32165) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(32165))))  severity failure;
	assert RAM(32166) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(32166))))  severity failure;
	assert RAM(32167) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(32167))))  severity failure;
	assert RAM(32168) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(32168))))  severity failure;
	assert RAM(32169) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(32169))))  severity failure;
	assert RAM(32170) = std_logic_vector(to_unsigned(23,8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(32170))))  severity failure;
	assert RAM(32171) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(32171))))  severity failure;
	assert RAM(32172) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(32172))))  severity failure;
	assert RAM(32173) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(32173))))  severity failure;
	assert RAM(32174) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(32174))))  severity failure;
	assert RAM(32175) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(32175))))  severity failure;
	assert RAM(32176) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(32176))))  severity failure;
	assert RAM(32177) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(32177))))  severity failure;
	assert RAM(32178) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(32178))))  severity failure;
	assert RAM(32179) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(32179))))  severity failure;
	assert RAM(32180) = std_logic_vector(to_unsigned(124,8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(32180))))  severity failure;
	assert RAM(32181) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(32181))))  severity failure;
	assert RAM(32182) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(32182))))  severity failure;
	assert RAM(32183) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(32183))))  severity failure;
	assert RAM(32184) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(32184))))  severity failure;
	assert RAM(32185) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(32185))))  severity failure;
	assert RAM(32186) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(32186))))  severity failure;
	assert RAM(32187) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(32187))))  severity failure;
	assert RAM(32188) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32188))))  severity failure;
	assert RAM(32189) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(32189))))  severity failure;
	assert RAM(32190) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(32190))))  severity failure;
	assert RAM(32191) = std_logic_vector(to_unsigned(65,8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(32191))))  severity failure;
	assert RAM(32192) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(32192))))  severity failure;
	assert RAM(32193) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(32193))))  severity failure;
	assert RAM(32194) = std_logic_vector(to_unsigned(131,8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(32194))))  severity failure;
	assert RAM(32195) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(32195))))  severity failure;
	assert RAM(32196) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(32196))))  severity failure;
	assert RAM(32197) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(32197))))  severity failure;
	assert RAM(32198) = std_logic_vector(to_unsigned(134,8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(32198))))  severity failure;
	assert RAM(32199) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(32199))))  severity failure;
	assert RAM(32200) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(32200))))  severity failure;
	assert RAM(32201) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(32201))))  severity failure;
	assert RAM(32202) = std_logic_vector(to_unsigned(176,8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(32202))))  severity failure;
	assert RAM(32203) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(32203))))  severity failure;
	assert RAM(32204) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(32204))))  severity failure;
	assert RAM(32205) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(32205))))  severity failure;
	assert RAM(32206) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(32206))))  severity failure;
	assert RAM(32207) = std_logic_vector(to_unsigned(177,8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(32207))))  severity failure;
	assert RAM(32208) = std_logic_vector(to_unsigned(110,8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(32208))))  severity failure;
	assert RAM(32209) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32209))))  severity failure;
	assert RAM(32210) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(32210))))  severity failure;
	assert RAM(32211) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(32211))))  severity failure;
	assert RAM(32212) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(32212))))  severity failure;
	assert RAM(32213) = std_logic_vector(to_unsigned(13,8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(32213))))  severity failure;
	assert RAM(32214) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(32214))))  severity failure;
	assert RAM(32215) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(32215))))  severity failure;
	assert RAM(32216) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(32216))))  severity failure;
	assert RAM(32217) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(32217))))  severity failure;
	assert RAM(32218) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32218))))  severity failure;
	assert RAM(32219) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(32219))))  severity failure;
	assert RAM(32220) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(32220))))  severity failure;
	assert RAM(32221) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(32221))))  severity failure;
	assert RAM(32222) = std_logic_vector(to_unsigned(58,8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(32222))))  severity failure;
	assert RAM(32223) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(32223))))  severity failure;
	assert RAM(32224) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(32224))))  severity failure;
	assert RAM(32225) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32225))))  severity failure;
	assert RAM(32226) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32226))))  severity failure;
	assert RAM(32227) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(32227))))  severity failure;
	assert RAM(32228) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(32228))))  severity failure;
	assert RAM(32229) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(32229))))  severity failure;
	assert RAM(32230) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32230))))  severity failure;
	assert RAM(32231) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32231))))  severity failure;
	assert RAM(32232) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(32232))))  severity failure;
	assert RAM(32233) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(32233))))  severity failure;
	assert RAM(32234) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(32234))))  severity failure;
	assert RAM(32235) = std_logic_vector(to_unsigned(118,8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(32235))))  severity failure;
	assert RAM(32236) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(32236))))  severity failure;
	assert RAM(32237) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(32237))))  severity failure;
	assert RAM(32238) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(32238))))  severity failure;
	assert RAM(32239) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32239))))  severity failure;
	assert RAM(32240) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(32240))))  severity failure;
	assert RAM(32241) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(32241))))  severity failure;
	assert RAM(32242) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(32242))))  severity failure;
	assert RAM(32243) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(32243))))  severity failure;
	assert RAM(32244) = std_logic_vector(to_unsigned(104,8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(32244))))  severity failure;
	assert RAM(32245) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32245))))  severity failure;
	assert RAM(32246) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(32246))))  severity failure;
	assert RAM(32247) = std_logic_vector(to_unsigned(218,8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(32247))))  severity failure;
	assert RAM(32248) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(32248))))  severity failure;
	assert RAM(32249) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(32249))))  severity failure;
	assert RAM(32250) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(32250))))  severity failure;
	assert RAM(32251) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(32251))))  severity failure;
	assert RAM(32252) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(32252))))  severity failure;
	assert RAM(32253) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(32253))))  severity failure;
	assert RAM(32254) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(32254))))  severity failure;
	assert RAM(32255) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(32255))))  severity failure;
	assert RAM(32256) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(32256))))  severity failure;
	assert RAM(32257) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32257))))  severity failure;
	assert RAM(32258) = std_logic_vector(to_unsigned(175,8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(32258))))  severity failure;
	assert RAM(32259) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32259))))  severity failure;
	assert RAM(32260) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32260))))  severity failure;
	assert RAM(32261) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(32261))))  severity failure;
	assert RAM(32262) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(32262))))  severity failure;
	assert RAM(32263) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(32263))))  severity failure;
	assert RAM(32264) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(32264))))  severity failure;
	assert RAM(32265) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(32265))))  severity failure;
	assert RAM(32266) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32266))))  severity failure;
	assert RAM(32267) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(32267))))  severity failure;
	assert RAM(32268) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(32268))))  severity failure;
	assert RAM(32269) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32269))))  severity failure;
	assert RAM(32270) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(32270))))  severity failure;
	assert RAM(32271) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(32271))))  severity failure;
	assert RAM(32272) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32272))))  severity failure;
	assert RAM(32273) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(32273))))  severity failure;
	assert RAM(32274) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(32274))))  severity failure;
	assert RAM(32275) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(32275))))  severity failure;
	assert RAM(32276) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(32276))))  severity failure;
	assert RAM(32277) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(32277))))  severity failure;
	assert RAM(32278) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(32278))))  severity failure;
	assert RAM(32279) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(32279))))  severity failure;
	assert RAM(32280) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(32280))))  severity failure;
	assert RAM(32281) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(32281))))  severity failure;
	assert RAM(32282) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32282))))  severity failure;
	assert RAM(32283) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(32283))))  severity failure;
	assert RAM(32284) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(32284))))  severity failure;
	assert RAM(32285) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(32285))))  severity failure;
	assert RAM(32286) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32286))))  severity failure;
	assert RAM(32287) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(32287))))  severity failure;
	assert RAM(32288) = std_logic_vector(to_unsigned(244,8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(32288))))  severity failure;
	assert RAM(32289) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(32289))))  severity failure;
	assert RAM(32290) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(32290))))  severity failure;
	assert RAM(32291) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(32291))))  severity failure;
	assert RAM(32292) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(32292))))  severity failure;
	assert RAM(32293) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(32293))))  severity failure;
	assert RAM(32294) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(32294))))  severity failure;
	assert RAM(32295) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(32295))))  severity failure;
	assert RAM(32296) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(32296))))  severity failure;
	assert RAM(32297) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(32297))))  severity failure;
	assert RAM(32298) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(32298))))  severity failure;
	assert RAM(32299) = std_logic_vector(to_unsigned(214,8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(32299))))  severity failure;
	assert RAM(32300) = std_logic_vector(to_unsigned(143,8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(32300))))  severity failure;
	assert RAM(32301) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(32301))))  severity failure;
	assert RAM(32302) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(32302))))  severity failure;
	assert RAM(32303) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32303))))  severity failure;
	assert RAM(32304) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32304))))  severity failure;
	assert RAM(32305) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(32305))))  severity failure;
	assert RAM(32306) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(32306))))  severity failure;
	assert RAM(32307) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(32307))))  severity failure;
	assert RAM(32308) = std_logic_vector(to_unsigned(99,8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(32308))))  severity failure;
	assert RAM(32309) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(32309))))  severity failure;
	assert RAM(32310) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(32310))))  severity failure;
	assert RAM(32311) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(32311))))  severity failure;
	assert RAM(32312) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(32312))))  severity failure;
	assert RAM(32313) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(32313))))  severity failure;
	assert RAM(32314) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(32314))))  severity failure;
	assert RAM(32315) = std_logic_vector(to_unsigned(112,8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(32315))))  severity failure;
	assert RAM(32316) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(32316))))  severity failure;
	assert RAM(32317) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(32317))))  severity failure;
	assert RAM(32318) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(32318))))  severity failure;
	assert RAM(32319) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(32319))))  severity failure;
	assert RAM(32320) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(32320))))  severity failure;
	assert RAM(32321) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(32321))))  severity failure;
	assert RAM(32322) = std_logic_vector(to_unsigned(84,8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(32322))))  severity failure;
	assert RAM(32323) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(32323))))  severity failure;
	assert RAM(32324) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(32324))))  severity failure;
	assert RAM(32325) = std_logic_vector(to_unsigned(15,8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(32325))))  severity failure;
	assert RAM(32326) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(32326))))  severity failure;
	assert RAM(32327) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(32327))))  severity failure;
	assert RAM(32328) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32328))))  severity failure;
	assert RAM(32329) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32329))))  severity failure;
	assert RAM(32330) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(32330))))  severity failure;
	assert RAM(32331) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(32331))))  severity failure;
	assert RAM(32332) = std_logic_vector(to_unsigned(106,8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(32332))))  severity failure;
	assert RAM(32333) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(32333))))  severity failure;
	assert RAM(32334) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32334))))  severity failure;
	assert RAM(32335) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(32335))))  severity failure;
	assert RAM(32336) = std_logic_vector(to_unsigned(116,8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(32336))))  severity failure;
	assert RAM(32337) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(32337))))  severity failure;
	assert RAM(32338) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(32338))))  severity failure;
	assert RAM(32339) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32339))))  severity failure;
	assert RAM(32340) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(32340))))  severity failure;
	assert RAM(32341) = std_logic_vector(to_unsigned(81,8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(32341))))  severity failure;
	assert RAM(32342) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(32342))))  severity failure;
	assert RAM(32343) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32343))))  severity failure;
	assert RAM(32344) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(32344))))  severity failure;
	assert RAM(32345) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(32345))))  severity failure;
	assert RAM(32346) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(32346))))  severity failure;
	assert RAM(32347) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32347))))  severity failure;
	assert RAM(32348) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(32348))))  severity failure;
	assert RAM(32349) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(32349))))  severity failure;
	assert RAM(32350) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32350))))  severity failure;
	assert RAM(32351) = std_logic_vector(to_unsigned(126,8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(32351))))  severity failure;
	assert RAM(32352) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(32352))))  severity failure;
	assert RAM(32353) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32353))))  severity failure;
	assert RAM(32354) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(32354))))  severity failure;
	assert RAM(32355) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(32355))))  severity failure;
	assert RAM(32356) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(32356))))  severity failure;
	assert RAM(32357) = std_logic_vector(to_unsigned(51,8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(32357))))  severity failure;
	assert RAM(32358) = std_logic_vector(to_unsigned(206,8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(32358))))  severity failure;
	assert RAM(32359) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(32359))))  severity failure;
	assert RAM(32360) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(32360))))  severity failure;
	assert RAM(32361) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32361))))  severity failure;
	assert RAM(32362) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(32362))))  severity failure;
	assert RAM(32363) = std_logic_vector(to_unsigned(45,8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(32363))))  severity failure;
	assert RAM(32364) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(32364))))  severity failure;
	assert RAM(32365) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(32365))))  severity failure;
	assert RAM(32366) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32366))))  severity failure;
	assert RAM(32367) = std_logic_vector(to_unsigned(36,8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(32367))))  severity failure;
	assert RAM(32368) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(32368))))  severity failure;
	assert RAM(32369) = std_logic_vector(to_unsigned(123,8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(32369))))  severity failure;
	assert RAM(32370) = std_logic_vector(to_unsigned(142,8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(32370))))  severity failure;
	assert RAM(32371) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(32371))))  severity failure;
	assert RAM(32372) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(32372))))  severity failure;
	assert RAM(32373) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(32373))))  severity failure;
	assert RAM(32374) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(32374))))  severity failure;
	assert RAM(32375) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(32375))))  severity failure;
	assert RAM(32376) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(32376))))  severity failure;
	assert RAM(32377) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(32377))))  severity failure;
	assert RAM(32378) = std_logic_vector(to_unsigned(238,8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(32378))))  severity failure;
	assert RAM(32379) = std_logic_vector(to_unsigned(174,8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(32379))))  severity failure;
	assert RAM(32380) = std_logic_vector(to_unsigned(156,8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(32380))))  severity failure;
	assert RAM(32381) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32381))))  severity failure;
	assert RAM(32382) = std_logic_vector(to_unsigned(119,8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(32382))))  severity failure;
	assert RAM(32383) = std_logic_vector(to_unsigned(31,8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(32383))))  severity failure;
	assert RAM(32384) = std_logic_vector(to_unsigned(187,8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(32384))))  severity failure;
	assert RAM(32385) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(32385))))  severity failure;
	assert RAM(32386) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32386))))  severity failure;
	assert RAM(32387) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(32387))))  severity failure;
	assert RAM(32388) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(32388))))  severity failure;
	assert RAM(32389) = std_logic_vector(to_unsigned(75,8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(32389))))  severity failure;
	assert RAM(32390) = std_logic_vector(to_unsigned(219,8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(32390))))  severity failure;
	assert RAM(32391) = std_logic_vector(to_unsigned(55,8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(32391))))  severity failure;
	assert RAM(32392) = std_logic_vector(to_unsigned(91,8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(32392))))  severity failure;
	assert RAM(32393) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32393))))  severity failure;
	assert RAM(32394) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(32394))))  severity failure;
	assert RAM(32395) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(32395))))  severity failure;
	assert RAM(32396) = std_logic_vector(to_unsigned(107,8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(32396))))  severity failure;
	assert RAM(32397) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(32397))))  severity failure;
	assert RAM(32398) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(32398))))  severity failure;
	assert RAM(32399) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(32399))))  severity failure;
	assert RAM(32400) = std_logic_vector(to_unsigned(146,8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(32400))))  severity failure;
	assert RAM(32401) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(32401))))  severity failure;
	assert RAM(32402) = std_logic_vector(to_unsigned(136,8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(32402))))  severity failure;
	assert RAM(32403) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(32403))))  severity failure;
	assert RAM(32404) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(32404))))  severity failure;
	assert RAM(32405) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(32405))))  severity failure;
	assert RAM(32406) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(32406))))  severity failure;
	assert RAM(32407) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(32407))))  severity failure;
	assert RAM(32408) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(32408))))  severity failure;
	assert RAM(32409) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32409))))  severity failure;
	assert RAM(32410) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32410))))  severity failure;
	assert RAM(32411) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(32411))))  severity failure;
	assert RAM(32412) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(32412))))  severity failure;
	assert RAM(32413) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(32413))))  severity failure;
	assert RAM(32414) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(32414))))  severity failure;
	assert RAM(32415) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(32415))))  severity failure;
	assert RAM(32416) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32416))))  severity failure;
	assert RAM(32417) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(32417))))  severity failure;
	assert RAM(32418) = std_logic_vector(to_unsigned(1,8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(32418))))  severity failure;
	assert RAM(32419) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(32419))))  severity failure;
	assert RAM(32420) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(32420))))  severity failure;
	assert RAM(32421) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32421))))  severity failure;
	assert RAM(32422) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(32422))))  severity failure;
	assert RAM(32423) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32423))))  severity failure;
	assert RAM(32424) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(32424))))  severity failure;
	assert RAM(32425) = std_logic_vector(to_unsigned(243,8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(32425))))  severity failure;
	assert RAM(32426) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(32426))))  severity failure;
	assert RAM(32427) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(32427))))  severity failure;
	assert RAM(32428) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(32428))))  severity failure;
	assert RAM(32429) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(32429))))  severity failure;
	assert RAM(32430) = std_logic_vector(to_unsigned(137,8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(32430))))  severity failure;
	assert RAM(32431) = std_logic_vector(to_unsigned(95,8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(32431))))  severity failure;
	assert RAM(32432) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(32432))))  severity failure;
	assert RAM(32433) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32433))))  severity failure;
	assert RAM(32434) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32434))))  severity failure;
	assert RAM(32435) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(32435))))  severity failure;
	assert RAM(32436) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32436))))  severity failure;
	assert RAM(32437) = std_logic_vector(to_unsigned(8,8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(32437))))  severity failure;
	assert RAM(32438) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(32438))))  severity failure;
	assert RAM(32439) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(32439))))  severity failure;
	assert RAM(32440) = std_logic_vector(to_unsigned(40,8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(32440))))  severity failure;
	assert RAM(32441) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(32441))))  severity failure;
	assert RAM(32442) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(32442))))  severity failure;
	assert RAM(32443) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(32443))))  severity failure;
	assert RAM(32444) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(32444))))  severity failure;
	assert RAM(32445) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(32445))))  severity failure;
	assert RAM(32446) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(32446))))  severity failure;
	assert RAM(32447) = std_logic_vector(to_unsigned(72,8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(32447))))  severity failure;
	assert RAM(32448) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32448))))  severity failure;
	assert RAM(32449) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(32449))))  severity failure;
	assert RAM(32450) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(32450))))  severity failure;
	assert RAM(32451) = std_logic_vector(to_unsigned(138,8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(32451))))  severity failure;
	assert RAM(32452) = std_logic_vector(to_unsigned(173,8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(32452))))  severity failure;
	assert RAM(32453) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(32453))))  severity failure;
	assert RAM(32454) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(32454))))  severity failure;
	assert RAM(32455) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32455))))  severity failure;
	assert RAM(32456) = std_logic_vector(to_unsigned(237,8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(32456))))  severity failure;
	assert RAM(32457) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(32457))))  severity failure;
	assert RAM(32458) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(32458))))  severity failure;
	assert RAM(32459) = std_logic_vector(to_unsigned(141,8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(32459))))  severity failure;
	assert RAM(32460) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(32460))))  severity failure;
	assert RAM(32461) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(32461))))  severity failure;
	assert RAM(32462) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32462))))  severity failure;
	assert RAM(32463) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(32463))))  severity failure;
	assert RAM(32464) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32464))))  severity failure;
	assert RAM(32465) = std_logic_vector(to_unsigned(102,8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(32465))))  severity failure;
	assert RAM(32466) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32466))))  severity failure;
	assert RAM(32467) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(32467))))  severity failure;
	assert RAM(32468) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(32468))))  severity failure;
	assert RAM(32469) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32469))))  severity failure;
	assert RAM(32470) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(32470))))  severity failure;
	assert RAM(32471) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(32471))))  severity failure;
	assert RAM(32472) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(32472))))  severity failure;
	assert RAM(32473) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(32473))))  severity failure;
	assert RAM(32474) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(32474))))  severity failure;
	assert RAM(32475) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(32475))))  severity failure;
	assert RAM(32476) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(32476))))  severity failure;
	assert RAM(32477) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(32477))))  severity failure;
	assert RAM(32478) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32478))))  severity failure;
	assert RAM(32479) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(32479))))  severity failure;
	assert RAM(32480) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(32480))))  severity failure;
	assert RAM(32481) = std_logic_vector(to_unsigned(19,8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(32481))))  severity failure;
	assert RAM(32482) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(32482))))  severity failure;
	assert RAM(32483) = std_logic_vector(to_unsigned(151,8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(32483))))  severity failure;
	assert RAM(32484) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(32484))))  severity failure;
	assert RAM(32485) = std_logic_vector(to_unsigned(215,8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(32485))))  severity failure;
	assert RAM(32486) = std_logic_vector(to_unsigned(209,8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(32486))))  severity failure;
	assert RAM(32487) = std_logic_vector(to_unsigned(222,8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(32487))))  severity failure;
	assert RAM(32488) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(32488))))  severity failure;
	assert RAM(32489) = std_logic_vector(to_unsigned(193,8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(32489))))  severity failure;
	assert RAM(32490) = std_logic_vector(to_unsigned(152,8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(32490))))  severity failure;
	assert RAM(32491) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(32491))))  severity failure;
	assert RAM(32492) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(32492))))  severity failure;
	assert RAM(32493) = std_logic_vector(to_unsigned(44,8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(32493))))  severity failure;
	assert RAM(32494) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(32494))))  severity failure;
	assert RAM(32495) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(32495))))  severity failure;
	assert RAM(32496) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(32496))))  severity failure;
	assert RAM(32497) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(32497))))  severity failure;
	assert RAM(32498) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(32498))))  severity failure;
	assert RAM(32499) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(32499))))  severity failure;
	assert RAM(32500) = std_logic_vector(to_unsigned(231,8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(32500))))  severity failure;
	assert RAM(32501) = std_logic_vector(to_unsigned(232,8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(32501))))  severity failure;
	assert RAM(32502) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(32502))))  severity failure;
	assert RAM(32503) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(32503))))  severity failure;
	assert RAM(32504) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(32504))))  severity failure;
	assert RAM(32505) = std_logic_vector(to_unsigned(108,8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(32505))))  severity failure;
	assert RAM(32506) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(32506))))  severity failure;
	assert RAM(32507) = std_logic_vector(to_unsigned(216,8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(32507))))  severity failure;
	assert RAM(32508) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32508))))  severity failure;
	assert RAM(32509) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(32509))))  severity failure;
	assert RAM(32510) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32510))))  severity failure;
	assert RAM(32511) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32511))))  severity failure;
	assert RAM(32512) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(32512))))  severity failure;
	assert RAM(32513) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32513))))  severity failure;
	assert RAM(32514) = std_logic_vector(to_unsigned(207,8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(32514))))  severity failure;
	assert RAM(32515) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(32515))))  severity failure;
	assert RAM(32516) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(32516))))  severity failure;
	assert RAM(32517) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(32517))))  severity failure;
	assert RAM(32518) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(32518))))  severity failure;
	assert RAM(32519) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(32519))))  severity failure;
	assert RAM(32520) = std_logic_vector(to_unsigned(194,8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(32520))))  severity failure;
	assert RAM(32521) = std_logic_vector(to_unsigned(111,8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(32521))))  severity failure;
	assert RAM(32522) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32522))))  severity failure;
	assert RAM(32523) = std_logic_vector(to_unsigned(12,8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(32523))))  severity failure;
	assert RAM(32524) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32524))))  severity failure;
	assert RAM(32525) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(32525))))  severity failure;
	assert RAM(32526) = std_logic_vector(to_unsigned(34,8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(32526))))  severity failure;
	assert RAM(32527) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(32527))))  severity failure;
	assert RAM(32528) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(32528))))  severity failure;
	assert RAM(32529) = std_logic_vector(to_unsigned(144,8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(32529))))  severity failure;
	assert RAM(32530) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(32530))))  severity failure;
	assert RAM(32531) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(32531))))  severity failure;
	assert RAM(32532) = std_logic_vector(to_unsigned(66,8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(32532))))  severity failure;
	assert RAM(32533) = std_logic_vector(to_unsigned(42,8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(32533))))  severity failure;
	assert RAM(32534) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(32534))))  severity failure;
	assert RAM(32535) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(32535))))  severity failure;
	assert RAM(32536) = std_logic_vector(to_unsigned(39,8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(32536))))  severity failure;
	assert RAM(32537) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(32537))))  severity failure;
	assert RAM(32538) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(32538))))  severity failure;
	assert RAM(32539) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32539))))  severity failure;
	assert RAM(32540) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32540))))  severity failure;
	assert RAM(32541) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(32541))))  severity failure;
	assert RAM(32542) = std_logic_vector(to_unsigned(52,8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(32542))))  severity failure;
	assert RAM(32543) = std_logic_vector(to_unsigned(127,8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(32543))))  severity failure;
	assert RAM(32544) = std_logic_vector(to_unsigned(189,8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(32544))))  severity failure;
	assert RAM(32545) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32545))))  severity failure;
	assert RAM(32546) = std_logic_vector(to_unsigned(247,8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(32546))))  severity failure;
	assert RAM(32547) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(32547))))  severity failure;
	assert RAM(32548) = std_logic_vector(to_unsigned(64,8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(32548))))  severity failure;
	assert RAM(32549) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(32549))))  severity failure;
	assert RAM(32550) = std_logic_vector(to_unsigned(183,8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(32550))))  severity failure;
	assert RAM(32551) = std_logic_vector(to_unsigned(109,8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(32551))))  severity failure;
	assert RAM(32552) = std_logic_vector(to_unsigned(97,8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(32552))))  severity failure;
	assert RAM(32553) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(32553))))  severity failure;
	assert RAM(32554) = std_logic_vector(to_unsigned(220,8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(32554))))  severity failure;
	assert RAM(32555) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32555))))  severity failure;
	assert RAM(32556) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(32556))))  severity failure;
	assert RAM(32557) = std_logic_vector(to_unsigned(70,8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(32557))))  severity failure;
	assert RAM(32558) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(32558))))  severity failure;
	assert RAM(32559) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(32559))))  severity failure;
	assert RAM(32560) = std_logic_vector(to_unsigned(87,8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(32560))))  severity failure;
	assert RAM(32561) = std_logic_vector(to_unsigned(249,8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(32561))))  severity failure;
	assert RAM(32562) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32562))))  severity failure;
	assert RAM(32563) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(32563))))  severity failure;
	assert RAM(32564) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(32564))))  severity failure;
	assert RAM(32565) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(32565))))  severity failure;
	assert RAM(32566) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(32566))))  severity failure;
	assert RAM(32567) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(32567))))  severity failure;
	assert RAM(32568) = std_logic_vector(to_unsigned(159,8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(32568))))  severity failure;
	assert RAM(32569) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(32569))))  severity failure;
	assert RAM(32570) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(32570))))  severity failure;
	assert RAM(32571) = std_logic_vector(to_unsigned(103,8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(32571))))  severity failure;
	assert RAM(32572) = std_logic_vector(to_unsigned(74,8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(32572))))  severity failure;
	assert RAM(32573) = std_logic_vector(to_unsigned(82,8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(32573))))  severity failure;
	assert RAM(32574) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(32574))))  severity failure;
	assert RAM(32575) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32575))))  severity failure;
	assert RAM(32576) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(32576))))  severity failure;
	assert RAM(32577) = std_logic_vector(to_unsigned(251,8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(32577))))  severity failure;
	assert RAM(32578) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32578))))  severity failure;
	assert RAM(32579) = std_logic_vector(to_unsigned(114,8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(32579))))  severity failure;
	assert RAM(32580) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(32580))))  severity failure;
	assert RAM(32581) = std_logic_vector(to_unsigned(154,8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(32581))))  severity failure;
	assert RAM(32582) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(32582))))  severity failure;
	assert RAM(32583) = std_logic_vector(to_unsigned(201,8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(32583))))  severity failure;
	assert RAM(32584) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(32584))))  severity failure;
	assert RAM(32585) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(32585))))  severity failure;
	assert RAM(32586) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(32586))))  severity failure;
	assert RAM(32587) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(32587))))  severity failure;
	assert RAM(32588) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(32588))))  severity failure;
	assert RAM(32589) = std_logic_vector(to_unsigned(17,8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(32589))))  severity failure;
	assert RAM(32590) = std_logic_vector(to_unsigned(213,8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(32590))))  severity failure;
	assert RAM(32591) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32591))))  severity failure;
	assert RAM(32592) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32592))))  severity failure;
	assert RAM(32593) = std_logic_vector(to_unsigned(24,8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(32593))))  severity failure;
	assert RAM(32594) = std_logic_vector(to_unsigned(43,8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(32594))))  severity failure;
	assert RAM(32595) = std_logic_vector(to_unsigned(205,8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(32595))))  severity failure;
	assert RAM(32596) = std_logic_vector(to_unsigned(85,8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(32596))))  severity failure;
	assert RAM(32597) = std_logic_vector(to_unsigned(16,8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(32597))))  severity failure;
	assert RAM(32598) = std_logic_vector(to_unsigned(182,8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(32598))))  severity failure;
	assert RAM(32599) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(32599))))  severity failure;
	assert RAM(32600) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(32600))))  severity failure;
	assert RAM(32601) = std_logic_vector(to_unsigned(133,8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(32601))))  severity failure;
	assert RAM(32602) = std_logic_vector(to_unsigned(241,8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(32602))))  severity failure;
	assert RAM(32603) = std_logic_vector(to_unsigned(128,8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(32603))))  severity failure;
	assert RAM(32604) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(32604))))  severity failure;
	assert RAM(32605) = std_logic_vector(to_unsigned(27,8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(32605))))  severity failure;
	assert RAM(32606) = std_logic_vector(to_unsigned(28,8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(32606))))  severity failure;
	assert RAM(32607) = std_logic_vector(to_unsigned(139,8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(32607))))  severity failure;
	assert RAM(32608) = std_logic_vector(to_unsigned(168,8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(32608))))  severity failure;
	assert RAM(32609) = std_logic_vector(to_unsigned(242,8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(32609))))  severity failure;
	assert RAM(32610) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32610))))  severity failure;
	assert RAM(32611) = std_logic_vector(to_unsigned(228,8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(32611))))  severity failure;
	assert RAM(32612) = std_logic_vector(to_unsigned(90,8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(32612))))  severity failure;
	assert RAM(32613) = std_logic_vector(to_unsigned(148,8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(32613))))  severity failure;
	assert RAM(32614) = std_logic_vector(to_unsigned(71,8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(32614))))  severity failure;
	assert RAM(32615) = std_logic_vector(to_unsigned(22,8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(32615))))  severity failure;
	assert RAM(32616) = std_logic_vector(to_unsigned(32,8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(32616))))  severity failure;
	assert RAM(32617) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32617))))  severity failure;
	assert RAM(32618) = std_logic_vector(to_unsigned(20,8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(32618))))  severity failure;
	assert RAM(32619) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32619))))  severity failure;
	assert RAM(32620) = std_logic_vector(to_unsigned(230,8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(32620))))  severity failure;
	assert RAM(32621) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(32621))))  severity failure;
	assert RAM(32622) = std_logic_vector(to_unsigned(0,8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(32622))))  severity failure;
	assert RAM(32623) = std_logic_vector(to_unsigned(120,8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(32623))))  severity failure;
	assert RAM(32624) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(32624))))  severity failure;
	assert RAM(32625) = std_logic_vector(to_unsigned(92,8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(32625))))  severity failure;
	assert RAM(32626) = std_logic_vector(to_unsigned(169,8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(32626))))  severity failure;
	assert RAM(32627) = std_logic_vector(to_unsigned(172,8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(32627))))  severity failure;
	assert RAM(32628) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(32628))))  severity failure;
	assert RAM(32629) = std_logic_vector(to_unsigned(252,8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(32629))))  severity failure;
	assert RAM(32630) = std_logic_vector(to_unsigned(6,8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(32630))))  severity failure;
	assert RAM(32631) = std_logic_vector(to_unsigned(100,8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(32631))))  severity failure;
	assert RAM(32632) = std_logic_vector(to_unsigned(96,8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(32632))))  severity failure;
	assert RAM(32633) = std_logic_vector(to_unsigned(224,8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(32633))))  severity failure;
	assert RAM(32634) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(32634))))  severity failure;
	assert RAM(32635) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32635))))  severity failure;
	assert RAM(32636) = std_logic_vector(to_unsigned(147,8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(32636))))  severity failure;
	assert RAM(32637) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(32637))))  severity failure;
	assert RAM(32638) = std_logic_vector(to_unsigned(165,8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(32638))))  severity failure;
	assert RAM(32639) = std_logic_vector(to_unsigned(61,8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(32639))))  severity failure;
	assert RAM(32640) = std_logic_vector(to_unsigned(76,8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(32640))))  severity failure;
	assert RAM(32641) = std_logic_vector(to_unsigned(83,8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(32641))))  severity failure;
	assert RAM(32642) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(32642))))  severity failure;
	assert RAM(32643) = std_logic_vector(to_unsigned(145,8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(32643))))  severity failure;
	assert RAM(32644) = std_logic_vector(to_unsigned(59,8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(32644))))  severity failure;
	assert RAM(32645) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32645))))  severity failure;
	assert RAM(32646) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32646))))  severity failure;
	assert RAM(32647) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32647))))  severity failure;
	assert RAM(32648) = std_logic_vector(to_unsigned(9,8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(32648))))  severity failure;
	assert RAM(32649) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32649))))  severity failure;
	assert RAM(32650) = std_logic_vector(to_unsigned(94,8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(32650))))  severity failure;
	assert RAM(32651) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32651))))  severity failure;
	assert RAM(32652) = std_logic_vector(to_unsigned(195,8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(32652))))  severity failure;
	assert RAM(32653) = std_logic_vector(to_unsigned(48,8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(32653))))  severity failure;
	assert RAM(32654) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(32654))))  severity failure;
	assert RAM(32655) = std_logic_vector(to_unsigned(73,8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(32655))))  severity failure;
	assert RAM(32656) = std_logic_vector(to_unsigned(190,8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(32656))))  severity failure;
	assert RAM(32657) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(32657))))  severity failure;
	assert RAM(32658) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(32658))))  severity failure;
	assert RAM(32659) = std_logic_vector(to_unsigned(86,8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(32659))))  severity failure;
	assert RAM(32660) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(32660))))  severity failure;
	assert RAM(32661) = std_logic_vector(to_unsigned(38,8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(32661))))  severity failure;
	assert RAM(32662) = std_logic_vector(to_unsigned(199,8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(32662))))  severity failure;
	assert RAM(32663) = std_logic_vector(to_unsigned(26,8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(32663))))  severity failure;
	assert RAM(32664) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(32664))))  severity failure;
	assert RAM(32665) = std_logic_vector(to_unsigned(135,8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(32665))))  severity failure;
	assert RAM(32666) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32666))))  severity failure;
	assert RAM(32667) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(32667))))  severity failure;
	assert RAM(32668) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(32668))))  severity failure;
	assert RAM(32669) = std_logic_vector(to_unsigned(226,8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(32669))))  severity failure;
	assert RAM(32670) = std_logic_vector(to_unsigned(121,8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(32670))))  severity failure;
	assert RAM(32671) = std_logic_vector(to_unsigned(253,8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(32671))))  severity failure;
	assert RAM(32672) = std_logic_vector(to_unsigned(132,8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(32672))))  severity failure;
	assert RAM(32673) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(32673))))  severity failure;
	assert RAM(32674) = std_logic_vector(to_unsigned(150,8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(32674))))  severity failure;
	assert RAM(32675) = std_logic_vector(to_unsigned(161,8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(32675))))  severity failure;
	assert RAM(32676) = std_logic_vector(to_unsigned(227,8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(32676))))  severity failure;
	assert RAM(32677) = std_logic_vector(to_unsigned(202,8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(32677))))  severity failure;
	assert RAM(32678) = std_logic_vector(to_unsigned(78,8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(32678))))  severity failure;
	assert RAM(32679) = std_logic_vector(to_unsigned(69,8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(32679))))  severity failure;
	assert RAM(32680) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32680))))  severity failure;
	assert RAM(32681) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32681))))  severity failure;
	assert RAM(32682) = std_logic_vector(to_unsigned(188,8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(32682))))  severity failure;
	assert RAM(32683) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(32683))))  severity failure;
	assert RAM(32684) = std_logic_vector(to_unsigned(57,8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(32684))))  severity failure;
	assert RAM(32685) = std_logic_vector(to_unsigned(250,8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(32685))))  severity failure;
	assert RAM(32686) = std_logic_vector(to_unsigned(210,8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(32686))))  severity failure;
	assert RAM(32687) = std_logic_vector(to_unsigned(37,8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(32687))))  severity failure;
	assert RAM(32688) = std_logic_vector(to_unsigned(117,8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(32688))))  severity failure;
	assert RAM(32689) = std_logic_vector(to_unsigned(35,8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(32689))))  severity failure;
	assert RAM(32690) = std_logic_vector(to_unsigned(60,8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(32690))))  severity failure;
	assert RAM(32691) = std_logic_vector(to_unsigned(80,8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(32691))))  severity failure;
	assert RAM(32692) = std_logic_vector(to_unsigned(255,8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(32692))))  severity failure;
	assert RAM(32693) = std_logic_vector(to_unsigned(50,8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(32693))))  severity failure;
	assert RAM(32694) = std_logic_vector(to_unsigned(192,8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(32694))))  severity failure;
	assert RAM(32695) = std_logic_vector(to_unsigned(89,8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(32695))))  severity failure;
	assert RAM(32696) = std_logic_vector(to_unsigned(245,8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(32696))))  severity failure;
	assert RAM(32697) = std_logic_vector(to_unsigned(93,8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(32697))))  severity failure;
	assert RAM(32698) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(32698))))  severity failure;
	assert RAM(32699) = std_logic_vector(to_unsigned(130,8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(32699))))  severity failure;
	assert RAM(32700) = std_logic_vector(to_unsigned(18,8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(32700))))  severity failure;
	assert RAM(32701) = std_logic_vector(to_unsigned(4,8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(32701))))  severity failure;
	assert RAM(32702) = std_logic_vector(to_unsigned(197,8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(32702))))  severity failure;
	assert RAM(32703) = std_logic_vector(to_unsigned(217,8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(32703))))  severity failure;
	assert RAM(32704) = std_logic_vector(to_unsigned(225,8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(32704))))  severity failure;
	assert RAM(32705) = std_logic_vector(to_unsigned(157,8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(32705))))  severity failure;
	assert RAM(32706) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(32706))))  severity failure;
	assert RAM(32707) = std_logic_vector(to_unsigned(11,8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(32707))))  severity failure;
	assert RAM(32708) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(32708))))  severity failure;
	assert RAM(32709) = std_logic_vector(to_unsigned(163,8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(32709))))  severity failure;
	assert RAM(32710) = std_logic_vector(to_unsigned(67,8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(32710))))  severity failure;
	assert RAM(32711) = std_logic_vector(to_unsigned(21,8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(32711))))  severity failure;
	assert RAM(32712) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32712))))  severity failure;
	assert RAM(32713) = std_logic_vector(to_unsigned(171,8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(32713))))  severity failure;
	assert RAM(32714) = std_logic_vector(to_unsigned(178,8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(32714))))  severity failure;
	assert RAM(32715) = std_logic_vector(to_unsigned(221,8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(32715))))  severity failure;
	assert RAM(32716) = std_logic_vector(to_unsigned(223,8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(32716))))  severity failure;
	assert RAM(32717) = std_logic_vector(to_unsigned(160,8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(32717))))  severity failure;
	assert RAM(32718) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(32718))))  severity failure;
	assert RAM(32719) = std_logic_vector(to_unsigned(47,8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(32719))))  severity failure;
	assert RAM(32720) = std_logic_vector(to_unsigned(164,8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(32720))))  severity failure;
	assert RAM(32721) = std_logic_vector(to_unsigned(180,8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(32721))))  severity failure;
	assert RAM(32722) = std_logic_vector(to_unsigned(185,8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(32722))))  severity failure;
	assert RAM(32723) = std_logic_vector(to_unsigned(166,8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(32723))))  severity failure;
	assert RAM(32724) = std_logic_vector(to_unsigned(211,8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(32724))))  severity failure;
	assert RAM(32725) = std_logic_vector(to_unsigned(41,8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(32725))))  severity failure;
	assert RAM(32726) = std_logic_vector(to_unsigned(140,8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(32726))))  severity failure;
	assert RAM(32727) = std_logic_vector(to_unsigned(10,8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(32727))))  severity failure;
	assert RAM(32728) = std_logic_vector(to_unsigned(181,8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(32728))))  severity failure;
	assert RAM(32729) = std_logic_vector(to_unsigned(7,8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(32729))))  severity failure;
	assert RAM(32730) = std_logic_vector(to_unsigned(54,8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(32730))))  severity failure;
	assert RAM(32731) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32731))))  severity failure;
	assert RAM(32732) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32732))))  severity failure;
	assert RAM(32733) = std_logic_vector(to_unsigned(179,8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(32733))))  severity failure;
	assert RAM(32734) = std_logic_vector(to_unsigned(30,8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(32734))))  severity failure;
	assert RAM(32735) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32735))))  severity failure;
	assert RAM(32736) = std_logic_vector(to_unsigned(149,8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(32736))))  severity failure;
	assert RAM(32737) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(32737))))  severity failure;
	assert RAM(32738) = std_logic_vector(to_unsigned(49,8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(32738))))  severity failure;
	assert RAM(32739) = std_logic_vector(to_unsigned(33,8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(32739))))  severity failure;
	assert RAM(32740) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(32740))))  severity failure;
	assert RAM(32741) = std_logic_vector(to_unsigned(68,8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(32741))))  severity failure;
	assert RAM(32742) = std_logic_vector(to_unsigned(79,8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(32742))))  severity failure;
	assert RAM(32743) = std_logic_vector(to_unsigned(186,8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(32743))))  severity failure;
	assert RAM(32744) = std_logic_vector(to_unsigned(101,8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(32744))))  severity failure;
	assert RAM(32745) = std_logic_vector(to_unsigned(239,8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(32745))))  severity failure;
	assert RAM(32746) = std_logic_vector(to_unsigned(63,8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(32746))))  severity failure;
	assert RAM(32747) = std_logic_vector(to_unsigned(246,8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(32747))))  severity failure;
	assert RAM(32748) = std_logic_vector(to_unsigned(46,8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(32748))))  severity failure;
	assert RAM(32749) = std_logic_vector(to_unsigned(129,8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(32749))))  severity failure;
	assert RAM(32750) = std_logic_vector(to_unsigned(212,8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(32750))))  severity failure;
	assert RAM(32751) = std_logic_vector(to_unsigned(236,8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(32751))))  severity failure;
	assert RAM(32752) = std_logic_vector(to_unsigned(208,8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(32752))))  severity failure;
	assert RAM(32753) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32753))))  severity failure;
	assert RAM(32754) = std_logic_vector(to_unsigned(191,8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(32754))))  severity failure;
	assert RAM(32755) = std_logic_vector(to_unsigned(248,8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(32755))))  severity failure;
	assert RAM(32756) = std_logic_vector(to_unsigned(234,8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(32756))))  severity failure;
	assert RAM(32757) = std_logic_vector(to_unsigned(113,8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(32757))))  severity failure;
	assert RAM(32758) = std_logic_vector(to_unsigned(122,8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(32758))))  severity failure;
	assert RAM(32759) = std_logic_vector(to_unsigned(203,8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(32759))))  severity failure;
	assert RAM(32760) = std_logic_vector(to_unsigned(233,8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(32760))))  severity failure;
	assert RAM(32761) = std_logic_vector(to_unsigned(53,8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(32761))))  severity failure;
	assert RAM(32762) = std_logic_vector(to_unsigned(196,8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(32762))))  severity failure;
	assert RAM(32763) = std_logic_vector(to_unsigned(2,8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(32763))))  severity failure;
	assert RAM(32764) = std_logic_vector(to_unsigned(162,8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(32764))))  severity failure;
	assert RAM(32765) = std_logic_vector(to_unsigned(167,8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(32765))))  severity failure;
	assert RAM(32766) = std_logic_vector(to_unsigned(229,8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(32766))))  severity failure;
	assert RAM(32767) = std_logic_vector(to_unsigned(29,8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(32767))))  severity failure;
	assert RAM(32768) = std_logic_vector(to_unsigned(235,8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(32768))))  severity failure;
	assert RAM(32769) = std_logic_vector(to_unsigned(105,8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(32769))))  severity failure;

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb; 


